
module fdiv(
    input wire [31:0] x1,
    input wire [31:0] x2,
    output wire [31:0] y);

    wire sa;
    wire [7:0] ea;
    wire [22:0] ma;
    assign sa = x2[31:31];
    assign ea = x2[30:23];
    assign ma = x2[22:0];

    wire [10:0] mal;
    assign mal = x2[22:12];

    wire [45:0] tdata;

    function [45:0] TDATA (
	input [10:0] MAL
    );
    begin
	casex(MAL)
        11'd0: TDATA = 46'b1111111111100000000000011111111110000000000001;
        11'd1: TDATA = 46'b1111111110100000000100111111111010000000011011;
        11'd2: TDATA = 46'b1111111101100000001100111111110110000001001011;
        11'd3: TDATA = 46'b1111111100100000011000011111110010000010010001;
        11'd4: TDATA = 46'b1111111011100000101000111111101110000011110011;
        11'd5: TDATA = 46'b1111111010100000111100011111101010000101101000;
        11'd6: TDATA = 46'b1111111001100001010100111111100110000111111010;
        11'd7: TDATA = 46'b1111111000100001110000111111100010001010100001;
        11'd8: TDATA = 46'b1111110111100010001111111111011110001101011101;
        11'd9: TDATA = 46'b1111110110100010110011111111011010010000110100;
        11'd10: TDATA = 46'b1111110101100011011100011111010110010100100100;
        11'd11: TDATA = 46'b1111110100100100000111111111010010011000101001;
        11'd12: TDATA = 46'b1111110011100100110111011111001110011101000101;
        11'd13: TDATA = 46'b1111110010100101101011011111001010100001111011;
        11'd14: TDATA = 46'b1111110001100110100001111111000110100111000011;
        11'd15: TDATA = 46'b1111110000100111011101011111000010101100100111;
        11'd16: TDATA = 46'b1111101111101000011100011110111110110010100000;
        11'd17: TDATA = 46'b1111101110101001011111011110111010111000110000;
        11'd18: TDATA = 46'b1111101101101010100111011110110110111111011101;
        11'd19: TDATA = 46'b1111101100101011110001111110110011000110011010;
        11'd20: TDATA = 46'b1111101011101101000000111110101111001101110010;
        11'd21: TDATA = 46'b1111101010101110010011011110101011010101011111;
        11'd22: TDATA = 46'b1111101001101111101001111110100111011101100011;
        11'd23: TDATA = 46'b1111101000110001000100011110100011100101111111;
        11'd24: TDATA = 46'b1111100111110010100011011110011111101110110101;
        11'd25: TDATA = 46'b1111100110110100000100111110011011110111111011;
        11'd26: TDATA = 46'b1111100101110101101010111110011000000001011100;
        11'd27: TDATA = 46'b1111100100110111010100011110010100001011010001;
        11'd28: TDATA = 46'b1111100011111001000011011110010000010101100100;
        11'd29: TDATA = 46'b1111100010111010110100011110001100100000000111;
        11'd30: TDATA = 46'b1111100001111100101001011110001000101011000001;
        11'd31: TDATA = 46'b1111100000111110100010111110000100110110010100;
        11'd32: TDATA = 46'b1111100000000000100000011110000001000001111110;
        11'd33: TDATA = 46'b1111011111000010100000011101111101001101111010;
        11'd34: TDATA = 46'b1111011110000100100101111101111001011010010011;
        11'd35: TDATA = 46'b1111011101000110101101111101110101100110111101;
        11'd36: TDATA = 46'b1111011100001000111001111101110001110011111110;
        11'd37: TDATA = 46'b1111011011001011001010111101101110000001011010;
        11'd38: TDATA = 46'b1111011010001101011101111101101010001111000110;
        11'd39: TDATA = 46'b1111011001001111110101111101100110011101001101;
        11'd40: TDATA = 46'b1111011000010010010000111101100010101011100111;
        11'd41: TDATA = 46'b1111010111010100110000011101011110111010011010;
        11'd42: TDATA = 46'b1111010110010111010011011101011011001001100010;
        11'd43: TDATA = 46'b1111010101011001111001111101010111011000111111;
        11'd44: TDATA = 46'b1111010100011100100100011101010011101000110100;
        11'd45: TDATA = 46'b1111010011011111010011011101001111111001000001;
        11'd46: TDATA = 46'b1111010010100010000100111101001100001001011111;
        11'd47: TDATA = 46'b1111010001100100111010111101001000011010010110;
        11'd48: TDATA = 46'b1111010000100111110011111101000100101011100001;
        11'd49: TDATA = 46'b1111001111101010110000111101000000111101000010;
        11'd50: TDATA = 46'b1111001110101101110010111100111101001110111110;
        11'd51: TDATA = 46'b1111001101110000110110111100111001100001001001;
        11'd52: TDATA = 46'b1111001100110011111111011100110101110011101101;
        11'd53: TDATA = 46'b1111001011110111001011111100110010000110100111;
        11'd54: TDATA = 46'b1111001010111010011010111100101110011001110011;
        11'd55: TDATA = 46'b1111001001111101101101111100101010101101010101;
        11'd56: TDATA = 46'b1111001001000001000101011100100111000001010001;
        11'd57: TDATA = 46'b1111001000000100100000011100100011010101100001;
        11'd58: TDATA = 46'b1111000111000111111111011100011111101010000111;
        11'd59: TDATA = 46'b1111000110001011100000111100011011111110111111;
        11'd60: TDATA = 46'b1111000101001111000110111100011000010100001111;
        11'd61: TDATA = 46'b1111000100010010110000011100010100101001110100;
        11'd62: TDATA = 46'b1111000011010110011101111100010000111111101111;
        11'd63: TDATA = 46'b1111000010011010001110111100001101010101111111;
        11'd64: TDATA = 46'b1111000001011110000011011100001001101100100100;
        11'd65: TDATA = 46'b1111000000100001111010111100000110000011011100;
        11'd66: TDATA = 46'b1110111111100101110110111100000010011010101100;
        11'd67: TDATA = 46'b1110111110101001110101111011111110110010001111;
        11'd68: TDATA = 46'b1110111101101101111000111011111011001010001000;
        11'd69: TDATA = 46'b1110111100110001111111111011110111100010011000;
        11'd70: TDATA = 46'b1110111011110110001001111011110011111010111010;
        11'd71: TDATA = 46'b1110111010111010010111111011110000010011110011;
        11'd72: TDATA = 46'b1110111001111110101001011011101100101101000000;
        11'd73: TDATA = 46'b1110111001000010111110111011101001000110100100;
        11'd74: TDATA = 46'b1110111000000111010110111011100101100000011000;
        11'd75: TDATA = 46'b1110110111001011110100011011100001111010101000;
        11'd76: TDATA = 46'b1110110110010000010011111011011110010101000111;
        11'd77: TDATA = 46'b1110110101010100110110111011011010101111111011;
        11'd78: TDATA = 46'b1110110100011001011101111011010111001011000101;
        11'd79: TDATA = 46'b1110110011011110001000011011010011100110100011;
        11'd80: TDATA = 46'b1110110010100010110111011011010000000010011001;
        11'd81: TDATA = 46'b1110110001100111101000011011001100011110011110;
        11'd82: TDATA = 46'b1110110000101100011101111011001000111010111011;
        11'd83: TDATA = 46'b1110101111110001010110111011000101010111101101;
        11'd84: TDATA = 46'b1110101110110110010010111011000001110100110000;
        11'd85: TDATA = 46'b1110101101111011010011011010111110010010001100;
        11'd86: TDATA = 46'b1110101101000000010110111010111010101111111010;
        11'd87: TDATA = 46'b1110101100000101011100111010110111001101111001;
        11'd88: TDATA = 46'b1110101011001010101000011010110011101100010011;
        11'd89: TDATA = 46'b1110101010001111110110111010110000001011000000;
        11'd90: TDATA = 46'b1110101001010101000111111010101100101001111101;
        11'd91: TDATA = 46'b1110101000011010011100011010101001001001001110;
        11'd92: TDATA = 46'b1110100111011111110101011010100101101000110111;
        11'd93: TDATA = 46'b1110100110100101010001011010100010001000110010;
        11'd94: TDATA = 46'b1110100101101010110000111010011110101001000001;
        11'd95: TDATA = 46'b1110100100110000010011111010011011001001100101;
        11'd96: TDATA = 46'b1110100011110101111010111010010111101010011110;
        11'd97: TDATA = 46'b1110100010111011100100011010010100001011101000;
        11'd98: TDATA = 46'b1110100010000001010011011010010000101101001101;
        11'd99: TDATA = 46'b1110100001000111000011111010001101001110111110;
        11'd100: TDATA = 46'b1110100000001100111000011010001001110001000110;
        11'd101: TDATA = 46'b1110011111010010101111111010000110010011011111;
        11'd102: TDATA = 46'b1110011110011000101011111010000010110110010000;
        11'd103: TDATA = 46'b1110011101011110101001111001111111011001010000;
        11'd104: TDATA = 46'b1110011100100100101100111001111011111100101001;
        11'd105: TDATA = 46'b1110011011101010110001111001111000100000010000;
        11'd106: TDATA = 46'b1110011010110000111011111001110101000100010000;
        11'd107: TDATA = 46'b1110011001110111000111111001110001101000011111;
        11'd108: TDATA = 46'b1110011000111101011000011001101110001101000110;
        11'd109: TDATA = 46'b1110011000000011101100011001101010110010000000;
        11'd110: TDATA = 46'b1110010111001010000010111001100111010111001010;
        11'd111: TDATA = 46'b1110010110010000011100111001100011111100101000;
        11'd112: TDATA = 46'b1110010101010110111011011001100000100010011110;
        11'd113: TDATA = 46'b1110010100011101011100011001011101001000100011;
        11'd114: TDATA = 46'b1110010011100100000000011001011001101110111011;
        11'd115: TDATA = 46'b1110010010101010101000111001010110010101101010;
        11'd116: TDATA = 46'b1110010001110001010100011001010010111100101010;
        11'd117: TDATA = 46'b1110010000111000000010111001001111100011111101;
        11'd118: TDATA = 46'b1110001111111110110100011001001100001011100001;
        11'd119: TDATA = 46'b1110001111000101101010111001001000110011011110;
        11'd120: TDATA = 46'b1110001110001100100010111001000101011011100111;
        11'd121: TDATA = 46'b1110001101010011100000011001000010000100001100;
        11'd122: TDATA = 46'b1110001100011010011111011000111110101100111101;
        11'd123: TDATA = 46'b1110001011100001100001111000111011010110000001;
        11'd124: TDATA = 46'b1110001010101000101000111000110111111111011100;
        11'd125: TDATA = 46'b1110001001101111110001011000110100101001000100;
        11'd126: TDATA = 46'b1110001000110110111111011000110001010011000110;
        11'd127: TDATA = 46'b1110000111111110001111011000101101111101010110;
        11'd128: TDATA = 46'b1110000111000101100011011000101010100111111100;
        11'd129: TDATA = 46'b1110000110001100111001111000100111010010110001;
        11'd130: TDATA = 46'b1110000101010100010100111000100011111101111110;
        11'd131: TDATA = 46'b1110000100011011110010111000100000101001011100;
        11'd132: TDATA = 46'b1110000011100011010011011000011101010101001010;
        11'd133: TDATA = 46'b1110000010101010110111011000011010000001001011;
        11'd134: TDATA = 46'b1110000001110010011111011000010110101101100001;
        11'd135: TDATA = 46'b1110000000111010001001111000010011011010000111;
        11'd136: TDATA = 46'b1110000000000001111000011000010000000111000010;
        11'd137: TDATA = 46'b1101111111001001101001111000001100110100001111;
        11'd138: TDATA = 46'b1101111110010001011110111000001001100001101110;
        11'd139: TDATA = 46'b1101111101011001010110111000000110001111011111;
        11'd140: TDATA = 46'b1101111100100001010001111000000010111101100010;
        11'd141: TDATA = 46'b1101111011101001010000110111111111101011111010;
        11'd142: TDATA = 46'b1101111010110001010010110111111100011010100011;
        11'd143: TDATA = 46'b1101111001111001011000010111111001001001011111;
        11'd144: TDATA = 46'b1101111001000001100000010111110101111000101011;
        11'd145: TDATA = 46'b1101111000001001101100010111110010101000001011;
        11'd146: TDATA = 46'b1101110111010001111011010111101111010111111101;
        11'd147: TDATA = 46'b1101110110011010001101010111101100001000000001;
        11'd148: TDATA = 46'b1101110101100010100011010111101000111000011001;
        11'd149: TDATA = 46'b1101110100101010111100010111100101101001000010;
        11'd150: TDATA = 46'b1101110011110011011000010111100010011001111101;
        11'd151: TDATA = 46'b1101110010111011110111010111011111001011001001;
        11'd152: TDATA = 46'b1101110010000100011001010111011011111100100110;
        11'd153: TDATA = 46'b1101110001001100111110110111011000101110010110;
        11'd154: TDATA = 46'b1101110000010101101000010111010101100000011011;
        11'd155: TDATA = 46'b1101101111011110010100010111010010010010101111;
        11'd156: TDATA = 46'b1101101110100111000011010111001111000101010101;
        11'd157: TDATA = 46'b1101101101101111110101010111001011111000001011;
        11'd158: TDATA = 46'b1101101100111000101011110111001000101011011001;
        11'd159: TDATA = 46'b1101101100000001100100110111000101011110110101;
        11'd160: TDATA = 46'b1101101011001010100000010111000010010010100001;
        11'd161: TDATA = 46'b1101101010010011100000010110111111000110100011;
        11'd162: TDATA = 46'b1101101001011100100010110110111011111010110100;
        11'd163: TDATA = 46'b1101101000100101101000010110111000101111010111;
        11'd164: TDATA = 46'b1101100111101110110000110110110101100100001010;
        11'd165: TDATA = 46'b1101100110110111111100110110110010011001010000;
        11'd166: TDATA = 46'b1101100110000001001100010110101111001110101001;
        11'd167: TDATA = 46'b1101100101001010011111010110101100000100010101;
        11'd168: TDATA = 46'b1101100100010011110100010110101000111010001110;
        11'd169: TDATA = 46'b1101100011011101001100110110100101110000011010;
        11'd170: TDATA = 46'b1101100010100110101000110110100010100110111000;
        11'd171: TDATA = 46'b1101100001110000000111110110011111011101101000;
        11'd172: TDATA = 46'b1101100000111001101001110110011100010100101000;
        11'd173: TDATA = 46'b1101100000000011001110110110011001001011111001;
        11'd174: TDATA = 46'b1101011111001100110111010110010110000011011101;
        11'd175: TDATA = 46'b1101011110010110100011010110010010111011010100;
        11'd176: TDATA = 46'b1101011101100000010001010110001111110011011000;
        11'd177: TDATA = 46'b1101011100101010000011010110001100101011110000;
        11'd178: TDATA = 46'b1101011011110011111000010110001001100100011001;
        11'd179: TDATA = 46'b1101011010111101101111110110000110011101010001;
        11'd180: TDATA = 46'b1101011010000111101010110110000011010110011011;
        11'd181: TDATA = 46'b1101011001010001101000110110000000001111110110;
        11'd182: TDATA = 46'b1101011000011011101010110101111101001001100110;
        11'd183: TDATA = 46'b1101010111100101101110110101111010000011100010;
        11'd184: TDATA = 46'b1101010110101111110101110101110110111101110000;
        11'd185: TDATA = 46'b1101010101111010000000110101110011111000010001;
        11'd186: TDATA = 46'b1101010101000100001111010101110000110011000110;
        11'd187: TDATA = 46'b1101010100001110011111010101101101101110000101;
        11'd188: TDATA = 46'b1101010011011000110011010101101010101001011000;
        11'd189: TDATA = 46'b1101010010100011001010110101100111100100111110;
        11'd190: TDATA = 46'b1101010001101101100100010101100100100000110001;
        11'd191: TDATA = 46'b1101010000111000000000110101100001011100110101;
        11'd192: TDATA = 46'b1101010000000010100000110101011110011001001011;
        11'd193: TDATA = 46'b1101001111001101000100110101011011010101110101;
        11'd194: TDATA = 46'b1101001110010111101010110101011000010010101100;
        11'd195: TDATA = 46'b1101001101100010010100010101010101001111110101;
        11'd196: TDATA = 46'b1101001100101100111111110101010010001101001100;
        11'd197: TDATA = 46'b1101001011110111101111010101001111001010110110;
        11'd198: TDATA = 46'b1101001011000010100001110101001100001000110001;
        11'd199: TDATA = 46'b1101001010001101010111010101001001000110111100;
        11'd200: TDATA = 46'b1101001001011000001111010101000110000101010110;
        11'd201: TDATA = 46'b1101001000100011001010110101000011000100000010;
        11'd202: TDATA = 46'b1101000111101110001000110101000000000010111101;
        11'd203: TDATA = 46'b1101000110111001001011010100111101000010001110;
        11'd204: TDATA = 46'b1101000110000100001111010100111010000001101010;
        11'd205: TDATA = 46'b1101000101001111010111010100110111000001011001;
        11'd206: TDATA = 46'b1101000100011010100001010100110100000001010110;
        11'd207: TDATA = 46'b1101000011100101101110110100110001000001100100;
        11'd208: TDATA = 46'b1101000010110000111111010100101110000010000011;
        11'd209: TDATA = 46'b1101000001111100010011010100101011000010110100;
        11'd210: TDATA = 46'b1101000001000111101001010100101000000011110010;
        11'd211: TDATA = 46'b1101000000010011000010110100100101000101000001;
        11'd212: TDATA = 46'b1100111111011110011101110100100010000110011100;
        11'd213: TDATA = 46'b1100111110101001111110110100011111001000010010;
        11'd214: TDATA = 46'b1100111101110101100000010100011100001010001111;
        11'd215: TDATA = 46'b1100111101000001000101110100011001001100100000;
        11'd216: TDATA = 46'b1100111100001100101101110100010110001110111111;
        11'd217: TDATA = 46'b1100111011011000011001010100010011010001110000;
        11'd218: TDATA = 46'b1100111010100100000111110100010000010100110001;
        11'd219: TDATA = 46'b1100111001101111111000110100001101011000000001;
        11'd220: TDATA = 46'b1100111000111011101100110100001010011011100001;
        11'd221: TDATA = 46'b1100111000000111100011110100000111011111010001;
        11'd222: TDATA = 46'b1100110111010011011101110100000100100011010001;
        11'd223: TDATA = 46'b1100110110011111011010110100000001100111100010;
        11'd224: TDATA = 46'b1100110101101011011011010011111110101100000100;
        11'd225: TDATA = 46'b1100110100110111011101110011111011110000110011;
        11'd226: TDATA = 46'b1100110100000011100011110011111000110101110011;
        11'd227: TDATA = 46'b1100110011001111101011110011110101111011000000;
        11'd228: TDATA = 46'b1100110010011011110111110011110011000000100001;
        11'd229: TDATA = 46'b1100110001101000000101010011110000000110001101;
        11'd230: TDATA = 46'b1100110000110100010111010011101101001100001101;
        11'd231: TDATA = 46'b1100110000000000101011010011101010010010011011;
        11'd232: TDATA = 46'b1100101111001101000010110011100111011000111010;
        11'd233: TDATA = 46'b1100101110011001011100110011100100011111100111;
        11'd234: TDATA = 46'b1100101101100101111001010011100001100110100010;
        11'd235: TDATA = 46'b1100101100110010011001010011011110101101101111;
        11'd236: TDATA = 46'b1100101011111110111100010011011011110101001100;
        11'd237: TDATA = 46'b1100101011001011100001110011011000111100110111;
        11'd238: TDATA = 46'b1100101010011000001010110011010110000100110100;
        11'd239: TDATA = 46'b1100101001100100110101110011010011001100111101;
        11'd240: TDATA = 46'b1100101000110001100011110011010000010101010110;
        11'd241: TDATA = 46'b1100100111111110010100110011001101011101111111;
        11'd242: TDATA = 46'b1100100111001011001000110011001010100110111000;
        11'd243: TDATA = 46'b1100100110010111111111110011000111110000000001;
        11'd244: TDATA = 46'b1100100101100100111001010011000100111001010111;
        11'd245: TDATA = 46'b1100100100110001110101010011000010000010111100;
        11'd246: TDATA = 46'b1100100011111110110100110010111111001100110010;
        11'd247: TDATA = 46'b1100100011001011110111110010111100010110111010;
        11'd248: TDATA = 46'b1100100010011000111100110010111001100001001110;
        11'd249: TDATA = 46'b1100100001100110000100110010110110101011110010;
        11'd250: TDATA = 46'b1100100000110011001111110010110011110110100110;
        11'd251: TDATA = 46'b1100100000000000011100110010110001000001100110;
        11'd252: TDATA = 46'b1100011111001101101101010010101110001100110111;
        11'd253: TDATA = 46'b1100011110011011000000010010101011011000010110;
        11'd254: TDATA = 46'b1100011101101000010110110010101000100100000111;
        11'd255: TDATA = 46'b1100011100110101101111010010100101110000000011;
        11'd256: TDATA = 46'b1100011100000011001011010010100010111100010010;
        11'd257: TDATA = 46'b1100011011010000101000110010100000001000101010;
        11'd258: TDATA = 46'b1100011010011110001011010010011101010101011001;
        11'd259: TDATA = 46'b1100011001101011101110110010011010100010010001;
        11'd260: TDATA = 46'b1100011000111001010101110010010111101111011010;
        11'd261: TDATA = 46'b1100011000000110111111010010010100111100110010;
        11'd262: TDATA = 46'b1100010111010100101011110010010010001010011000;
        11'd263: TDATA = 46'b1100010110100010011011010010001111011000001110;
        11'd264: TDATA = 46'b1100010101110000001100110010001100100110010001;
        11'd265: TDATA = 46'b1100010100111110000010110010001001110100101000;
        11'd266: TDATA = 46'b1100010100001011111001010010000111000011000101;
        11'd267: TDATA = 46'b1100010011011001110011110010000100010001110110;
        11'd268: TDATA = 46'b1100010010100111110000110010000001100000110101;
        11'd269: TDATA = 46'b1100010001110101110000010001111110110000000001;
        11'd270: TDATA = 46'b1100010001000011110011010001111011111111011111;
        11'd271: TDATA = 46'b1100010000010001111000110001111001001111001010;
        11'd272: TDATA = 46'b1100001111100000000000110001110110011111000011;
        11'd273: TDATA = 46'b1100001110101110001100010001110011101111001101;
        11'd274: TDATA = 46'b1100001101111100011001010001110000111111100001;
        11'd275: TDATA = 46'b1100001101001010101001010001101110010000000101;
        11'd276: TDATA = 46'b1100001100011000111100010001101011100000111000;
        11'd277: TDATA = 46'b1100001011100111010010110001101000110001111100;
        11'd278: TDATA = 46'b1100001010110101101011010001100110000011001100;
        11'd279: TDATA = 46'b1100001010000100000101110001100011010100101000;
        11'd280: TDATA = 46'b1100001001010010100100010001100000100110010111;
        11'd281: TDATA = 46'b1100001000100001000100110001011101111000010010;
        11'd282: TDATA = 46'b1100000111101111101001010001011011001010011111;
        11'd283: TDATA = 46'b1100000110111110001110110001011000011100110101;
        11'd284: TDATA = 46'b1100000110001100111000010001010101101111011110;
        11'd285: TDATA = 46'b1100000101011011100011110001010011000010010010;
        11'd286: TDATA = 46'b1100000100101010010001110001010000010101010100;
        11'd287: TDATA = 46'b1100000011111001000010110001001101101000100101;
        11'd288: TDATA = 46'b1100000011000111110111010001001010111100001000;
        11'd289: TDATA = 46'b1100000010010110101100110001001000001111110010;
        11'd290: TDATA = 46'b1100000001100101100101110001000101100011101101;
        11'd291: TDATA = 46'b1100000000110100100001110001000010110111111000;
        11'd292: TDATA = 46'b1100000000000011100000010001000000001100010000;
        11'd293: TDATA = 46'b1011111111010010100001110000111101100000110111;
        11'd294: TDATA = 46'b1011111110100001100101010000111010110101101010;
        11'd295: TDATA = 46'b1011111101110000101011110000111000001010101100;
        11'd296: TDATA = 46'b1011111100111111110100110000110101011111111100;
        11'd297: TDATA = 46'b1011111100001111000000010000110010110101011001;
        11'd298: TDATA = 46'b1011111011011110001111010000110000001011000110;
        11'd299: TDATA = 46'b1011111010101101100000110000101101100001000010;
        11'd300: TDATA = 46'b1011111001111100110100010000101010110111001000;
        11'd301: TDATA = 46'b1011111001001100001010110000101000001101011110;
        11'd302: TDATA = 46'b1011111000011011100100010000100101100100000011;
        11'd303: TDATA = 46'b1011110111101011000000010000100010111010110101;
        11'd304: TDATA = 46'b1011110110111010011101110000100000010001110010;
        11'd305: TDATA = 46'b1011110110001001111111010000011101101001000000;
        11'd306: TDATA = 46'b1011110101011001100010110000011011000000011010;
        11'd307: TDATA = 46'b1011110100101001001000110000011000011000000010;
        11'd308: TDATA = 46'b1011110011111000110001110000010101101111111000;
        11'd309: TDATA = 46'b1011110011001000011101110000010011000111111110;
        11'd310: TDATA = 46'b1011110010011000001011110000010000100000001111;
        11'd311: TDATA = 46'b1011110001100111111100110000001101111000101110;
        11'd312: TDATA = 46'b1011110000110111110000010000001011010001011100;
        11'd313: TDATA = 46'b1011110000000111100110110000001000101010011000;
        11'd314: TDATA = 46'b1011101111010111011110110000000110000011011101;
        11'd315: TDATA = 46'b1011101110100111011001110000000011011100110010;
        11'd316: TDATA = 46'b1011101101110111011000010000000000110110010111;
        11'd317: TDATA = 46'b1011101101000111011000001111111110010000000111;
        11'd318: TDATA = 46'b1011101100010111011011001111111011101010000100;
        11'd319: TDATA = 46'b1011101011100111100000101111111001000100010000;
        11'd320: TDATA = 46'b1011101010110111101001001111110110011110101010;
        11'd321: TDATA = 46'b1011101010000111110100001111110011111001010001;
        11'd322: TDATA = 46'b1011101001011000000001001111110001010100000011;
        11'd323: TDATA = 46'b1011101000101000010001001111101110101111000100;
        11'd324: TDATA = 46'b1011100111111000100100001111101100001010010100;
        11'd325: TDATA = 46'b1011100111001000111000101111101001100101101110;
        11'd326: TDATA = 46'b1011100110011001010000001111100111000001010111;
        11'd327: TDATA = 46'b1011100101101001101010101111100100011101001110;
        11'd328: TDATA = 46'b1011100100111010001000001111100001111001010100;
        11'd329: TDATA = 46'b1011100100001010100111101111011111010101100101;
        11'd330: TDATA = 46'b1011100011011011001000001111011100110001111110;
        11'd331: TDATA = 46'b1011100010101011101101001111011010001110101011;
        11'd332: TDATA = 46'b1011100001111100010100101111010111101011100110;
        11'd333: TDATA = 46'b1011100001001100111101101111010101001000101001;
        11'd334: TDATA = 46'b1011100000011101101001101111010010100101111100;
        11'd335: TDATA = 46'b1011011111101110011000101111010000000011011101;
        11'd336: TDATA = 46'b1011011110111111001001101111001101100001001001;
        11'd337: TDATA = 46'b1011011110001111111101101111001010111111000100;
        11'd338: TDATA = 46'b1011011101100000110100101111001000011101001101;
        11'd339: TDATA = 46'b1011011100110001101101001111000101111011100000;
        11'd340: TDATA = 46'b1011011100000010101000001111000011011010000000;
        11'd341: TDATA = 46'b1011011011010011100111001111000000111000110010;
        11'd342: TDATA = 46'b1011011010100100100111001110111110010111101100;
        11'd343: TDATA = 46'b1011011001110101101001001110111011110110110001;
        11'd344: TDATA = 46'b1011011001000110101110101110111001010110000110;
        11'd345: TDATA = 46'b1011011000010111110111001110110110110101101010;
        11'd346: TDATA = 46'b1011010111101001000001001110110100010101010111;
        11'd347: TDATA = 46'b1011010110111010001101101110110001110101010001;
        11'd348: TDATA = 46'b1011010110001011011101001110101111010101011001;
        11'd349: TDATA = 46'b1011010101011100101111101110101100110101110001;
        11'd350: TDATA = 46'b1011010100101110000100001110101010010110010011;
        11'd351: TDATA = 46'b1011010011111111011010101110100111110111000000;
        11'd352: TDATA = 46'b1011010011010000110100101110100101010111111101;
        11'd353: TDATA = 46'b1011010010100010010000001110100010111001000100;
        11'd354: TDATA = 46'b1011010001110011101101101110100000011010010110;
        11'd355: TDATA = 46'b1011010001000101001111101110011101111011111011;
        11'd356: TDATA = 46'b1011010000010110110010101110011011011101101001;
        11'd357: TDATA = 46'b1011001111101000011000001110011000111111100010;
        11'd358: TDATA = 46'b1011001110111010000000101110010110100001101010;
        11'd359: TDATA = 46'b1011001110001011101011001110010100000011111110;
        11'd360: TDATA = 46'b1011001101011101011000001110010001100110011110;
        11'd361: TDATA = 46'b1011001100101111001000001110001111001001001100;
        11'd362: TDATA = 46'b1011001100000000111001101110001100101100000011;
        11'd363: TDATA = 46'b1011001011010010101111001110001010001111001101;
        11'd364: TDATA = 46'b1011001010100100100101101110000111110010011110;
        11'd365: TDATA = 46'b1011001001110110011110101110000101010101111011;
        11'd366: TDATA = 46'b1011001001001000011010101110000010111001100111;
        11'd367: TDATA = 46'b1011001000011010011000101110000000011101011110;
        11'd368: TDATA = 46'b1011000111101100011010101101111110000001100110;
        11'd369: TDATA = 46'b1011000110111110011100101101111011100101110011;
        11'd370: TDATA = 46'b1011000110010000100010101101111001001010010001;
        11'd371: TDATA = 46'b1011000101100010101010101101110110101110111010;
        11'd372: TDATA = 46'b1011000100110100110101001101110100010011110000;
        11'd373: TDATA = 46'b1011000100000111000001101101110001111000110001;
        11'd374: TDATA = 46'b1011000011011001010001001101101111011101111111;
        11'd375: TDATA = 46'b1011000010101011100011001101101101000011011011;
        11'd376: TDATA = 46'b1011000001111101110111101101101010101001000011;
        11'd377: TDATA = 46'b1011000001010000001110101101101000001110110111;
        11'd378: TDATA = 46'b1011000000100010100110101101100101110100110011;
        11'd379: TDATA = 46'b1010111111110101000001101101100011011010111101;
        11'd380: TDATA = 46'b1010111111000111100000001101100001000001010111;
        11'd381: TDATA = 46'b1010111110011010000000001101011110100111111010;
        11'd382: TDATA = 46'b1010111101101100100010101101011100001110101010;
        11'd383: TDATA = 46'b1010111100111111001000001101011001110101100111;
        11'd384: TDATA = 46'b1010111100010001101111101101010111011100110000;
        11'd385: TDATA = 46'b1010111011100100011000101101010101000100000001;
        11'd386: TDATA = 46'b1010111010110111000100101101010010101011100001;
        11'd387: TDATA = 46'b1010111010001001110011101101010000010011001111;
        11'd388: TDATA = 46'b1010111001011100100100101101001101111011000111;
        11'd389: TDATA = 46'b1010111000101111011000001101001011100011001100;
        11'd390: TDATA = 46'b1010111000000010001101101101001001001011011011;
        11'd391: TDATA = 46'b1010110111010101000101001101000110110011110110;
        11'd392: TDATA = 46'b1010110110101000000000001101000100011100100000;
        11'd393: TDATA = 46'b1010110101111010111100101101000010000101010011;
        11'd394: TDATA = 46'b1010110101001101111011101100111111101110010010;
        11'd395: TDATA = 46'b1010110100100000111100101100111101010111011100;
        11'd396: TDATA = 46'b1010110011110100000000101100111011000000110100;
        11'd397: TDATA = 46'b1010110011000111000110101100111000101010010110;
        11'd398: TDATA = 46'b1010110010011010001111101100110110010100000111;
        11'd399: TDATA = 46'b1010110001101101011010101100110011111110000010;
        11'd400: TDATA = 46'b1010110001000000100111101100110001101000001000;
        11'd401: TDATA = 46'b1010110000010011110111001100101111010010011010;
        11'd402: TDATA = 46'b1010101111100111001000101100101100111100110111;
        11'd403: TDATA = 46'b1010101110111010011101001100101010100111100010;
        11'd404: TDATA = 46'b1010101110001101110011101100101000010010010111;
        11'd405: TDATA = 46'b1010101101100001001100101100100101111101011000;
        11'd406: TDATA = 46'b1010101100110100101000001100100011101000100110;
        11'd407: TDATA = 46'b1010101100001000000101001100100001010011111101;
        11'd408: TDATA = 46'b1010101011011011100100101100011110111111100000;
        11'd409: TDATA = 46'b1010101010101111000111001100011100101011010000;
        11'd410: TDATA = 46'b1010101010000010101011101100011010010111001011;
        11'd411: TDATA = 46'b1010101001010110010010101100011000000011010011;
        11'd412: TDATA = 46'b1010101000101001111100001100010101101111100110;
        11'd413: TDATA = 46'b1010100111111101100111001100010011011100000011;
        11'd414: TDATA = 46'b1010100111010001010101001100010001001000101101;
        11'd415: TDATA = 46'b1010100110100101000100101100001110110101100000;
        11'd416: TDATA = 46'b1010100101111000110111001100001100100010100001;
        11'd417: TDATA = 46'b1010100101001100101100001100001010001111101110;
        11'd418: TDATA = 46'b1010100100100000100010101100000111111101000100;
        11'd419: TDATA = 46'b1010100011110100011100001100000101101010100111;
        11'd420: TDATA = 46'b1010100011001000011000001100000011011000010111;
        11'd421: TDATA = 46'b1010100010011100010100101100000001000110001100;
        11'd422: TDATA = 46'b1010100001110000010100101011111110110100010000;
        11'd423: TDATA = 46'b1010100001000100010111101011111100100010100010;
        11'd424: TDATA = 46'b1010100000011000011011101011111010010000111100;
        11'd425: TDATA = 46'b1010011111101100100010101011110111111111100011;
        11'd426: TDATA = 46'b1010011111000000101100001011110101101110010110;
        11'd427: TDATA = 46'b1010011110010100110111101011110011011101010011;
        11'd428: TDATA = 46'b1010011101101001000101001011110001001100011011;
        11'd429: TDATA = 46'b1010011100111101010101001011101110111011101111;
        11'd430: TDATA = 46'b1010011100010001100111001011101100101011001101;
        11'd431: TDATA = 46'b1010011011100101111100001011101010011010111000;
        11'd432: TDATA = 46'b1010011010111010010010101011101000001010101101;
        11'd433: TDATA = 46'b1010011010001110101011001011100101111010101100;
        11'd434: TDATA = 46'b1010011001100011000110101011100011101010111000;
        11'd435: TDATA = 46'b1010011000110111100100001011100001011011001111;
        11'd436: TDATA = 46'b1010011000001100000011101011011111001011110000;
        11'd437: TDATA = 46'b1010010111100000100110101011011100111100100000;
        11'd438: TDATA = 46'b1010010110110101001001101011011010101101010100;
        11'd439: TDATA = 46'b1010010110001001110000001011011000011110010111;
        11'd440: TDATA = 46'b1010010101011110011000101011010110001111100100;
        11'd441: TDATA = 46'b1010010100110011000100001011010100000000111111;
        11'd442: TDATA = 46'b1010010100000111110001001011010001110010100011;
        11'd443: TDATA = 46'b1010010011011100100000001011001111100100010000;
        11'd444: TDATA = 46'b1010010010110001010001101011001101010110001010;
        11'd445: TDATA = 46'b1010010010000110000101001011001011001000001110;
        11'd446: TDATA = 46'b1010010001011010111011101011001000111010011111;
        11'd447: TDATA = 46'b1010010000101111110011101011000110101100111001;
        11'd448: TDATA = 46'b1010010000000100101101101011000100011111011101;
        11'd449: TDATA = 46'b1010001111011001101010101011000010010010001111;
        11'd450: TDATA = 46'b1010001110101110101001001011000000000101001001;
        11'd451: TDATA = 46'b1010001110000011101011001010111101111000010010;
        11'd452: TDATA = 46'b1010001101011000101101101010111011101011100001;
        11'd453: TDATA = 46'b1010001100101101110011001010111001011110111100;
        11'd454: TDATA = 46'b1010001100000010111010101010110111010010100011;
        11'd455: TDATA = 46'b1010001011011000000100101010110101000110010100;
        11'd456: TDATA = 46'b1010001010101101010000001010110010111010001111;
        11'd457: TDATA = 46'b1010001010000010011111001010110000101110011000;
        11'd458: TDATA = 46'b1010001001010111101111001010101110100010101000;
        11'd459: TDATA = 46'b1010001000101101000001101010101100010111000100;
        11'd460: TDATA = 46'b1010001000000010010110101010101010001011101011;
        11'd461: TDATA = 46'b1010000111010111101101101010101000000000011101;
        11'd462: TDATA = 46'b1010000110101101000110101010100101110101011001;
        11'd463: TDATA = 46'b1010000110000010100001101010100011101010011111;
        11'd464: TDATA = 46'b1010000101010111111111101010100001011111110010;
        11'd465: TDATA = 46'b1010000100101101011111001010011111010101001110;
        11'd466: TDATA = 46'b1010000100000011000000001010011101001010110010;
        11'd467: TDATA = 46'b1010000011011000100100101010011011000000100100;
        11'd468: TDATA = 46'b1010000010101110001010101010011000110110100000;
        11'd469: TDATA = 46'b1010000010000011110010101010010110101100100101;
        11'd470: TDATA = 46'b1010000001011001011101001010010100100010110110;
        11'd471: TDATA = 46'b1010000000101111001001101010010010011001010001;
        11'd472: TDATA = 46'b1010000000000100111000001010010000001111110110;
        11'd473: TDATA = 46'b1001111111011010101001001010001110000110100111;
        11'd474: TDATA = 46'b1001111110110000011100001010001011111101100001;
        11'd475: TDATA = 46'b1001111110000110010001001010001001110100100110;
        11'd476: TDATA = 46'b1001111101011100001000001010000111101011110100;
        11'd477: TDATA = 46'b1001111100110010000001101010000101100011001110;
        11'd478: TDATA = 46'b1001111100000111111101001010000011011010110010;
        11'd479: TDATA = 46'b1001111011011101111011001010000001010010100010;
        11'd480: TDATA = 46'b1001111010110011111011001001111111001010011011;
        11'd481: TDATA = 46'b1001111010001001111100001001111101000010011100;
        11'd482: TDATA = 46'b1001111001100000000000101001111010111010101011;
        11'd483: TDATA = 46'b1001111000110110000110101001111000110011000010;
        11'd484: TDATA = 46'b1001111000001100001111001001110110101011100101;
        11'd485: TDATA = 46'b1001110111100010011001001001110100100100010000;
        11'd486: TDATA = 46'b1001110110111000100101101001110010011101000110;
        11'd487: TDATA = 46'b1001110110001110110100101001110000010110001000;
        11'd488: TDATA = 46'b1001110101100101000101001001101110001111010011;
        11'd489: TDATA = 46'b1001110100111011011000001001101100001000101000;
        11'd490: TDATA = 46'b1001110100010001101100101001101010000010000110;
        11'd491: TDATA = 46'b1001110011101000000100001001100111111011110001;
        11'd492: TDATA = 46'b1001110010111110011101001001100101110101100101;
        11'd493: TDATA = 46'b1001110010010100111000001001100011101111100010;
        11'd494: TDATA = 46'b1001110001101011010101001001100001101001101001;
        11'd495: TDATA = 46'b1001110001000001110100101001011111100011111011;
        11'd496: TDATA = 46'b1001110000011000010110101001011101011110011001;
        11'd497: TDATA = 46'b1001101111101110111001101001011011011000111101;
        11'd498: TDATA = 46'b1001101111000101100000001001011001010011110000;
        11'd499: TDATA = 46'b1001101110011100000111101001010111001110101010;
        11'd500: TDATA = 46'b1001101101110010110001001001010101001001101101;
        11'd501: TDATA = 46'b1001101101001001011101101001010011000100111101;
        11'd502: TDATA = 46'b1001101100100000001011001001010001000000010100;
        11'd503: TDATA = 46'b1001101011110110111011001001001110111011110111;
        11'd504: TDATA = 46'b1001101011001101101100101001001100110111100001;
        11'd505: TDATA = 46'b1001101010100100100001001001001010110011011000;
        11'd506: TDATA = 46'b1001101001111011010111101001001000101111011001;
        11'd507: TDATA = 46'b1001101001010010001111101001000110101011100010;
        11'd508: TDATA = 46'b1001101000101001001001101001000100100111110101;
        11'd509: TDATA = 46'b1001101000000000000110101001000010100100010101;
        11'd510: TDATA = 46'b1001100111010111000100101001000000100000111011;
        11'd511: TDATA = 46'b1001100110101110000101101000111110011101101110;
        11'd512: TDATA = 46'b1001100110000101001000001000111100011010101001;
        11'd513: TDATA = 46'b1001100101011100001100101000111010010111101110;
        11'd514: TDATA = 46'b1001100100110011010011101000111000010100111110;
        11'd515: TDATA = 46'b1001100100001010011100001000110110010010010111;
        11'd516: TDATA = 46'b1001100011100001100111001000110100001111111010;
        11'd517: TDATA = 46'b1001100010111000110011101000110010001101100110;
        11'd518: TDATA = 46'b1001100010010000000010101000110000001011011100;
        11'd519: TDATA = 46'b1001100001100111010011101000101110001001011101;
        11'd520: TDATA = 46'b1001100000111110100101101000101100000111100011;
        11'd521: TDATA = 46'b1001100000010101111011101000101010000101111010;
        11'd522: TDATA = 46'b1001011111101101010001101000101000000100010100;
        11'd523: TDATA = 46'b1001011111000100101010101000100110000010111011;
        11'd524: TDATA = 46'b1001011110011100000101101000100100000001101011;
        11'd525: TDATA = 46'b1001011101110011100010101000100010000000100101;
        11'd526: TDATA = 46'b1001011101001011000001001000011111111111100111;
        11'd527: TDATA = 46'b1001011100100010100011001000011101111110110111;
        11'd528: TDATA = 46'b1001011011111010000101101000011011111110001101;
        11'd529: TDATA = 46'b1001011011010001101010101000011001111101101101;
        11'd530: TDATA = 46'b1001011010101001010001101000010111111101010110;
        11'd531: TDATA = 46'b1001011010000000111011001000010101111101001011;
        11'd532: TDATA = 46'b1001011001011000100110101000010011111101001010;
        11'd533: TDATA = 46'b1001011000110000010011001000010001111101001111;
        11'd534: TDATA = 46'b1001011000001000000001101000001111111101011101;
        11'd535: TDATA = 46'b1001010111011111110011101000001101111101111001;
        11'd536: TDATA = 46'b1001010110110111100101101000001011111110011001;
        11'd537: TDATA = 46'b1001010110001111011011101000001001111111001001;
        11'd538: TDATA = 46'b1001010101100111010010101000000111111111111110;
        11'd539: TDATA = 46'b1001010100111111001011001000000110000000111100;
        11'd540: TDATA = 46'b1001010100010111000101101000000100000010000011;
        11'd541: TDATA = 46'b1001010011101111000011101000000010000011011001;
        11'd542: TDATA = 46'b1001010011000111000010101000000000000100110101;
        11'd543: TDATA = 46'b1001010010011111000011000111111110000110011000;
        11'd544: TDATA = 46'b1001010001110111000101100111111100001000000101;
        11'd545: TDATA = 46'b1001010001001111001010100111111010001001111101;
        11'd546: TDATA = 46'b1001010000100111010001000111111000001011111101;
        11'd547: TDATA = 46'b1001001111111111011010100111110110001110001010;
        11'd548: TDATA = 46'b1001001111010111100100100111110100010000011011;
        11'd549: TDATA = 46'b1001001110101111110001100111110010010010111001;
        11'd550: TDATA = 46'b1001001110001000000000100111110000010101100000;
        11'd551: TDATA = 46'b1001001101100000010001000111101110011000001111;
        11'd552: TDATA = 46'b1001001100111000100100000111101100011011001000;
        11'd553: TDATA = 46'b1001001100010000111000000111101010011110001001;
        11'd554: TDATA = 46'b1001001011101001001111000111101000100001010101;
        11'd555: TDATA = 46'b1001001011000001100111000111100110100100101000;
        11'd556: TDATA = 46'b1001001010011010000001100111100100101000000110;
        11'd557: TDATA = 46'b1001001001110010011101100111100010101011101011;
        11'd558: TDATA = 46'b1001001001001010111100000111100000101111011100;
        11'd559: TDATA = 46'b1001001000100011011100000111011110110011010100;
        11'd560: TDATA = 46'b1001000111111011111111000111011100110111011001;
        11'd561: TDATA = 46'b1001000111010100100010100111011010111011100010;
        11'd562: TDATA = 46'b1001000110101101001000100111011000111111110110;
        11'd563: TDATA = 46'b1001000110000101110000100111010111000100010100;
        11'd564: TDATA = 46'b1001000101011110011011000111010101001000111100;
        11'd565: TDATA = 46'b1001000100110111000110100111010011001101101011;
        11'd566: TDATA = 46'b1001000100001111110100000111010001010010100011;
        11'd567: TDATA = 46'b1001000011101000100011100111001111010111100100;
        11'd568: TDATA = 46'b1001000011000001010101100111001101011100110000;
        11'd569: TDATA = 46'b1001000010011010001000100111001011100010000010;
        11'd570: TDATA = 46'b1001000001110010111110100111001001100111100000;
        11'd571: TDATA = 46'b1001000001001011110101100111000111101101000101;
        11'd572: TDATA = 46'b1001000000100100101111000111000101110010110100;
        11'd573: TDATA = 46'b1000111111111101101001100111000011111000101010;
        11'd574: TDATA = 46'b1000111111010110101000000111000001111110101111;
        11'd575: TDATA = 46'b1000111110101111100101100111000000000100110100;
        11'd576: TDATA = 46'b1000111110001000100111100110111110001011001001;
        11'd577: TDATA = 46'b1000111101100001101010100110111100010001100101;
        11'd578: TDATA = 46'b1000111100111010101110100110111010011000000111;
        11'd579: TDATA = 46'b1000111100010011110101000110111000011110110100;
        11'd580: TDATA = 46'b1000111011101100111101000110110110100101101001;
        11'd581: TDATA = 46'b1000111011000110001000000110110100101100101001;
        11'd582: TDATA = 46'b1000111010011111010100000110110010110011110000;
        11'd583: TDATA = 46'b1000111001111000100010100110110000111011000001;
        11'd584: TDATA = 46'b1000111001010001110010100110101111000010011011;
        11'd585: TDATA = 46'b1000111000101011000100000110101101001001111011;
        11'd586: TDATA = 46'b1000111000000100011000000110101011010001100111;
        11'd587: TDATA = 46'b1000110111011101101101100110101001011001011010;
        11'd588: TDATA = 46'b1000110110110111000101000110100111100001010110;
        11'd589: TDATA = 46'b1000110110010000011110100110100101101001011011;
        11'd590: TDATA = 46'b1000110101101001111001100110100011110001101000;
        11'd591: TDATA = 46'b1000110101000011010111100110100001111010000001;
        11'd592: TDATA = 46'b1000110100011100110101100110100000000010011101;
        11'd593: TDATA = 46'b1000110011110110010111100110011110001011001000;
        11'd594: TDATA = 46'b1000110011001111111001100110011100010011110110;
        11'd595: TDATA = 46'b1000110010101001011110100110011010011100110000;
        11'd596: TDATA = 46'b1000110010000011000100100110011000100101110001;
        11'd597: TDATA = 46'b1000110001011100101100100110010110101110111010;
        11'd598: TDATA = 46'b1000110000110110010111000110010100111000001110;
        11'd599: TDATA = 46'b1000110000010000000011100110010011000001101011;
        11'd600: TDATA = 46'b1000101111101001110001100110010001001011010000;
        11'd601: TDATA = 46'b1000101111000011100001000110001111010100111100;
        11'd602: TDATA = 46'b1000101110011101010010100110001101011110110001;
        11'd603: TDATA = 46'b1000101101110111000101100110001011101000101101;
        11'd604: TDATA = 46'b1000101101010000111011100110001001110010110110;
        11'd605: TDATA = 46'b1000101100101010110011000110000111111101000110;
        11'd606: TDATA = 46'b1000101100000100101011100110000110000111011100;
        11'd607: TDATA = 46'b1000101011011110100110100110000100010001111101;
        11'd608: TDATA = 46'b1000101010111000100011100110000010011100100111;
        11'd609: TDATA = 46'b1000101010010010100001000110000000100111010101;
        11'd610: TDATA = 46'b1000101001101100100001000101111110110010001101;
        11'd611: TDATA = 46'b1000101001000110100100000101111100111101010010;
        11'd612: TDATA = 46'b1000101000100000100111100101111011001000011011;
        11'd613: TDATA = 46'b1000100111111010101101100101111001010011101110;
        11'd614: TDATA = 46'b1000100111010100110100100101110111011111000111;
        11'd615: TDATA = 46'b1000100110101110111111000101110101101010101110;
        11'd616: TDATA = 46'b1000100110001001001001100101110011110110011000;
        11'd617: TDATA = 46'b1000100101100011010111000101110010000010001110;
        11'd618: TDATA = 46'b1000100100111101100101100101110000001110001001;
        11'd619: TDATA = 46'b1000100100010111110110100101101110011010001111;
        11'd620: TDATA = 46'b1000100011110010001000100101101100100110011011;
        11'd621: TDATA = 46'b1000100011001100011101000101101010110010110010;
        11'd622: TDATA = 46'b1000100010100110110011100101101000111111010001;
        11'd623: TDATA = 46'b1000100010000001001011100101100111001011111000;
        11'd624: TDATA = 46'b1000100001011011100101000101100101011000100110;
        11'd625: TDATA = 46'b1000100000110110000000100101100011100101011100;
        11'd626: TDATA = 46'b1000100000010000011101100101100001110010011011;
        11'd627: TDATA = 46'b1000011111101010111100100101011111111111100010;
        11'd628: TDATA = 46'b1000011111000101011110100101011110001100110101;
        11'd629: TDATA = 46'b1000011110100000000000000101011100011010001001;
        11'd630: TDATA = 46'b1000011101111010100101000101011010100111101011;
        11'd631: TDATA = 46'b1000011101010101001011100101011000110101010100;
        11'd632: TDATA = 46'b1000011100101111110011100101010111000011000100;
        11'd633: TDATA = 46'b1000011100001010011101000101010101010000111100;
        11'd634: TDATA = 46'b1000011011100101001000000101010011011110111011;
        11'd635: TDATA = 46'b1000011010111111110110100101010001101101000111;
        11'd636: TDATA = 46'b1000011010011010100101100101001111111011011000;
        11'd637: TDATA = 46'b1000011001110101010110100101001110001001110001;
        11'd638: TDATA = 46'b1000011001010000001000100101001100011000010000;
        11'd639: TDATA = 46'b1000011000101010111101000101001010100110111010;
        11'd640: TDATA = 46'b1000011000000101110011100101001000110101101100;
        11'd641: TDATA = 46'b1000010111100000101011100101000111000100100101;
        11'd642: TDATA = 46'b1000010110111011100101100101000101010011101000;
        11'd643: TDATA = 46'b1000010110010110100001000101000011100010110001;
        11'd644: TDATA = 46'b1000010101110001011111000101000001110010000101;
        11'd645: TDATA = 46'b1000010101001100011101000101000000000001011100;
        11'd646: TDATA = 46'b1000010100100111011110100100111110010001000000;
        11'd647: TDATA = 46'b1000010100000010100001000100111100100000101001;
        11'd648: TDATA = 46'b1000010011011101100101100100111010110000011100;
        11'd649: TDATA = 46'b1000010010111000101100000100111001000000010111;
        11'd650: TDATA = 46'b1000010010010011110011100100110111010000010111;
        11'd651: TDATA = 46'b1000010001101110111100100100110101100000011111;
        11'd652: TDATA = 46'b1000010001001010001000000100110011110000110010;
        11'd653: TDATA = 46'b1000010000100101010101100100110010000001001101;
        11'd654: TDATA = 46'b1000010000000000100100100100110000010001101111;
        11'd655: TDATA = 46'b1000001111011011110101000100101110100010011000;
        11'd656: TDATA = 46'b1000001110110111001000000100101100110011001011;
        11'd657: TDATA = 46'b1000001110010010011100000100101011000100000101;
        11'd658: TDATA = 46'b1000001101101101110001000100101001010101000011;
        11'd659: TDATA = 46'b1000001101001001001001000100100111100110001110;
        11'd660: TDATA = 46'b1000001100100100100010100100100101110111100000;
        11'd661: TDATA = 46'b1000001011111111111101000100100100001000110111;
        11'd662: TDATA = 46'b1000001011011011011001100100100010011010010111;
        11'd663: TDATA = 46'b1000001010110110111000100100100000101100000001;
        11'd664: TDATA = 46'b1000001010010010011000000100011110111101101111;
        11'd665: TDATA = 46'b1000001001101101111010100100011101001111101001;
        11'd666: TDATA = 46'b1000001001001001011110100100011011100001101010;
        11'd667: TDATA = 46'b1000001000100101000011000100011001110011101111;
        11'd668: TDATA = 46'b1000001000000000101001100100011000000101111101;
        11'd669: TDATA = 46'b1000000111011100010011000100010110011000010111;
        11'd670: TDATA = 46'b1000000110110111111101100100010100101010110110;
        11'd671: TDATA = 46'b1000000110010011101010100100010010111101011111;
        11'd672: TDATA = 46'b1000000101101111010111100100010001010000001010;
        11'd673: TDATA = 46'b1000000101001011000111000100001111100011000000;
        11'd674: TDATA = 46'b1000000100100110111000100100001101110101111110;
        11'd675: TDATA = 46'b1000000100000010101100000100001100001001000101;
        11'd676: TDATA = 46'b1000000011011110100000000100001010011100010000;
        11'd677: TDATA = 46'b1000000010111010010111000100001000101111100111;
        11'd678: TDATA = 46'b1000000010010110001111000100000111000011000011;
        11'd679: TDATA = 46'b1000000001110010001000100100000101010110100110;
        11'd680: TDATA = 46'b1000000001001110000100000100000011101010010010;
        11'd681: TDATA = 46'b1000000000101010000001000100000001111110000101;
        11'd682: TDATA = 46'b1000000000000110000000000100000000010010000000;
        11'd683: TDATA = 46'b0111111111100010000000000011111110100110000001;
        11'd684: TDATA = 46'b0111111110111110000011000011111100111010001101;
        11'd685: TDATA = 46'b0111111110011010000111000011111011001110011111;
        11'd686: TDATA = 46'b0111111101110110001100100011111001100010111000;
        11'd687: TDATA = 46'b0111111101010010010011100011110111110111011000;
        11'd688: TDATA = 46'b0111111100101110011100100011110110001100000000;
        11'd689: TDATA = 46'b0111111100001010100111100011110100100000110001;
        11'd690: TDATA = 46'b0111111011100110110100000011110010110101101001;
        11'd691: TDATA = 46'b0111111011000011000001100011110001001010100111;
        11'd692: TDATA = 46'b0111111010011111010001100011101111011111101110;
        11'd693: TDATA = 46'b0111111001111011100010100011101101110100111011;
        11'd694: TDATA = 46'b0111111001010111110101100011101100001010010000;
        11'd695: TDATA = 46'b0111111000110100001011000011101010011111101111;
        11'd696: TDATA = 46'b0111111000010000100000100011101000110101010001;
        11'd697: TDATA = 46'b0111110111101100111001000011100111001010111110;
        11'd698: TDATA = 46'b0111110111001001010010100011100101100000110001;
        11'd699: TDATA = 46'b0111110110100101101101100011100011110110101011;
        11'd700: TDATA = 46'b0111110110000010001010100011100010001100101101;
        11'd701: TDATA = 46'b0111110101011110101000100011100000100010110100;
        11'd702: TDATA = 46'b0111110100111011001010100011011110111001001010;
        11'd703: TDATA = 46'b0111110100010111101011100011011101001111100000;
        11'd704: TDATA = 46'b0111110011110100001111000011011011100101111111;
        11'd705: TDATA = 46'b0111110011010000110100000011011001111100100101;
        11'd706: TDATA = 46'b0111110010101101011011100011011000010011010101;
        11'd707: TDATA = 46'b0111110010001010000100000011010110101010001010;
        11'd708: TDATA = 46'b0111110001100110101101100011010101000001000101;
        11'd709: TDATA = 46'b0111110001000011011001100011010011011000001010;
        11'd710: TDATA = 46'b0111110000100000000111100011010001101111010111;
        11'd711: TDATA = 46'b0111101111111100110101100011010000000110100111;
        11'd712: TDATA = 46'b0111101111011001100111000011001110011110000011;
        11'd713: TDATA = 46'b0111101110110110011000100011001100110101100010;
        11'd714: TDATA = 46'b0111101110010011001101000011001011001101001100;
        11'd715: TDATA = 46'b0111101101110000000011100011001001100100111111;
        11'd716: TDATA = 46'b0111101101001100111010100011000111111100110101;
        11'd717: TDATA = 46'b0111101100101001110011000011000110010100110010;
        11'd718: TDATA = 46'b0111101100000110101101100011000100101100111000;
        11'd719: TDATA = 46'b0111101011100011101001100011000011000101000100;
        11'd720: TDATA = 46'b0111101011000000101000000011000001011101011010;
        11'd721: TDATA = 46'b0111101010011101100111000010111111110101110100;
        11'd722: TDATA = 46'b0111101001111010101000000010111110001110010111;
        11'd723: TDATA = 46'b0111101001010111101010100010111100100111000000;
        11'd724: TDATA = 46'b0111101000110100101110100010111010111111110000;
        11'd725: TDATA = 46'b0111101000010001110100100010111001011000101000;
        11'd726: TDATA = 46'b0111100111101110111011100010110111110001100110;
        11'd727: TDATA = 46'b0111100111001100000100100010110110001010101100;
        11'd728: TDATA = 46'b0111100110101001001111100010110100100011111010;
        11'd729: TDATA = 46'b0111100110000110011011100010110010111101001110;
        11'd730: TDATA = 46'b0111100101100011101001100010110001010110101001;
        11'd731: TDATA = 46'b0111100101000000111000100010101111110000001011;
        11'd732: TDATA = 46'b0111100100011110001001100010101110001001110100;
        11'd733: TDATA = 46'b0111100011111011011100000010101100100011100100;
        11'd734: TDATA = 46'b0111100011011000110000100010101010111101011100;
        11'd735: TDATA = 46'b0111100010110110000111000010101001010111011101;
        11'd736: TDATA = 46'b0111100010010011011110100010100111110001100011;
        11'd737: TDATA = 46'b0111100001110000110111000010100110001011101110;
        11'd738: TDATA = 46'b0111100001001110010001100010100100100110000001;
        11'd739: TDATA = 46'b0111100000101011101101100010100011000000011100;
        11'd740: TDATA = 46'b0111100000001001001100000010100001011010111111;
        11'd741: TDATA = 46'b0111011111100110101011100010011111110101101000;
        11'd742: TDATA = 46'b0111011111000100001100000010011110010000010111;
        11'd743: TDATA = 46'b0111011110100001101110100010011100101011001101;
        11'd744: TDATA = 46'b0111011101111111010010100010011011000110001011;
        11'd745: TDATA = 46'b0111011101011100111000000010011001100001001110;
        11'd746: TDATA = 46'b0111011100111010011111100010010111111100011011;
        11'd747: TDATA = 46'b0111011100011000001000100010010110010111101101;
        11'd748: TDATA = 46'b0111011011110101110011000010010100110011000111;
        11'd749: TDATA = 46'b0111011011010011011111000010010011001110100111;
        11'd750: TDATA = 46'b0111011010110001001100100010010001101010001110;
        11'd751: TDATA = 46'b0111011010001110111011100010010000000101111100;
        11'd752: TDATA = 46'b0111011001101100101100100010001110100001110010;
        11'd753: TDATA = 46'b0111011001001010011110100010001100111101101101;
        11'd754: TDATA = 46'b0111011000101000010010100010001011011001110000;
        11'd755: TDATA = 46'b0111011000000110001000000010001001110101111001;
        11'd756: TDATA = 46'b0111010111100011111111000010001000010010001010;
        11'd757: TDATA = 46'b0111010111000001110111000010000110101110011111;
        11'd758: TDATA = 46'b0111010110011111110001000010000101001010111101;
        11'd759: TDATA = 46'b0111010101111101101100100010000011100111100010;
        11'd760: TDATA = 46'b0111010101011011101001100010000010000100001101;
        11'd761: TDATA = 46'b0111010100111001101000100010000000100001000000;
        11'd762: TDATA = 46'b0111010100010111101000100001111110111101111000;
        11'd763: TDATA = 46'b0111010011110101101011000001111101011010111010;
        11'd764: TDATA = 46'b0111010011010011101110100001111011111000000001;
        11'd765: TDATA = 46'b0111010010110001110011000001111010010101001101;
        11'd766: TDATA = 46'b0111010010001111111001000001111000110010100000;
        11'd767: TDATA = 46'b0111010001101110000001000001110111001111111011;
        11'd768: TDATA = 46'b0111010001001100001011000001110101101101011110;
        11'd769: TDATA = 46'b0111010000101010010110100001110100001011000111;
        11'd770: TDATA = 46'b0111010000001000100010100001110010101000110100;
        11'd771: TDATA = 46'b0111001111100110110000000001110001000110101000;
        11'd772: TDATA = 46'b0111001111000101000000100001101111100100100111;
        11'd773: TDATA = 46'b0111001110100011010001100001101110000010101001;
        11'd774: TDATA = 46'b0111001110000001100100000001101100100000110010;
        11'd775: TDATA = 46'b0111001101011111111000000001101010111111000010;
        11'd776: TDATA = 46'b0111001100111110001110100001101001011101011011;
        11'd777: TDATA = 46'b0111001100011100100101100001100111111011110111;
        11'd778: TDATA = 46'b0111001011111010111110100001100110011010011100;
        11'd779: TDATA = 46'b0111001011011001011000100001100100111001000110;
        11'd780: TDATA = 46'b0111001010110111110100100001100011010111111000;
        11'd781: TDATA = 46'b0111001010010110010001100001100001110110101111;
        11'd782: TDATA = 46'b0111001001110100110000100001100000010101101110;
        11'd783: TDATA = 46'b0111001001010011010001000001011110110100110011;
        11'd784: TDATA = 46'b0111001000110001110011100001011101010100000000;
        11'd785: TDATA = 46'b0111001000010000010110100001011011110011010001;
        11'd786: TDATA = 46'b0111000111101110111011100001011010010010101010;
        11'd787: TDATA = 46'b0111000111001101100001100001011000110010001000;
        11'd788: TDATA = 46'b0111000110101100001001100001010111010001101110;
        11'd789: TDATA = 46'b0111000110001010110011100001010101110001011100;
        11'd790: TDATA = 46'b0111000101101001011111000001010100010001010001;
        11'd791: TDATA = 46'b0111000101001000001011100001010010110001001010;
        11'd792: TDATA = 46'b0111000100100110111001000001010001010001001001;
        11'd793: TDATA = 46'b0111000100000101101000100001001111110001001111;
        11'd794: TDATA = 46'b0111000011100100011001100001001110010001011100;
        11'd795: TDATA = 46'b0111000011000011001100000001001100110001110000;
        11'd796: TDATA = 46'b0111000010100010000000000001001011010010001010;
        11'd797: TDATA = 46'b0111000010000000110101000001001001110010101001;
        11'd798: TDATA = 46'b0111000001011111101100100001001000010011010001;
        11'd799: TDATA = 46'b0111000000111110100100100001000110110011111101;
        11'd800: TDATA = 46'b0111000000011101011110100001000101010100110001;
        11'd801: TDATA = 46'b0110111111111100011001100001000011110101101001;
        11'd802: TDATA = 46'b0110111111011011010111000001000010010110101011;
        11'd803: TDATA = 46'b0110111110111010010101000001000000110111110001;
        11'd804: TDATA = 46'b0110111110011001010101000000111111011000111111;
        11'd805: TDATA = 46'b0110111101111000010111000000111101111010010100;
        11'd806: TDATA = 46'b0110111101010111011001100000111100011011101101;
        11'd807: TDATA = 46'b0110111100110110011101100000111010111101001100;
        11'd808: TDATA = 46'b0110111100010101100011100000111001011110110100;
        11'd809: TDATA = 46'b0110111011110100101010100000111000000000100000;
        11'd810: TDATA = 46'b0110111011010011110011100000110110100010010100;
        11'd811: TDATA = 46'b0110111010110010111101100000110101000100001101;
        11'd812: TDATA = 46'b0110111010010010001001000000110011100110001101;
        11'd813: TDATA = 46'b0110111001110001010110100000110010001000010100;
        11'd814: TDATA = 46'b0110111001010000100101000000110000101010100000;
        11'd815: TDATA = 46'b0110111000101111110101000000101111001100110011;
        11'd816: TDATA = 46'b0110111000001111000110100000101101101111001100;
        11'd817: TDATA = 46'b0110110111101110011001100000101100010001101011;
        11'd818: TDATA = 46'b0110110111001101101101100000101010110100010000;
        11'd819: TDATA = 46'b0110110110101101000100000000101001010110111101;
        11'd820: TDATA = 46'b0110110110001100011011100000100111111001110000;
        11'd821: TDATA = 46'b0110110101101011110100100000100110011100101001;
        11'd822: TDATA = 46'b0110110101001011001110100000100100111111100110;
        11'd823: TDATA = 46'b0110110100101010101001100000100011100010101001;
        11'd824: TDATA = 46'b0110110100001010001000000000100010000101111000;
        11'd825: TDATA = 46'b0110110011101001100101100000100000101001000110;
        11'd826: TDATA = 46'b0110110011001001000110100000011111001100100000;
        11'd827: TDATA = 46'b0110110010101000100111100000011101101111111100;
        11'd828: TDATA = 46'b0110110010001000001010100000011100010011100000;
        11'd829: TDATA = 46'b0110110001100111101111000000011010110111001010;
        11'd830: TDATA = 46'b0110110001000111010101000000011001011010111011;
        11'd831: TDATA = 46'b0110110000100110111100000000010111111110110000;
        11'd832: TDATA = 46'b0110110000000110100100100000010110100010101100;
        11'd833: TDATA = 46'b0110101111100110001111000000010101000110101111;
        11'd834: TDATA = 46'b0110101111000101111011000000010011101010111001;
        11'd835: TDATA = 46'b0110101110100101100111100000010010001111000110;
        11'd836: TDATA = 46'b0110101110000101010110100000010000110011011101;
        11'd837: TDATA = 46'b0110101101100101000110100000001111010111111000;
        11'd838: TDATA = 46'b0110101101000100110111100000001101111100011000;
        11'd839: TDATA = 46'b0110101100100100101001100000001100100000111101;
        11'd840: TDATA = 46'b0110101100000100011111000000001011000101101110;
        11'd841: TDATA = 46'b0110101011100100010100000000001001101010011111;
        11'd842: TDATA = 46'b0110101011000100001011100000001000001111011010;
        11'd843: TDATA = 46'b0110101010100100000011100000000110110100011000;
        11'd844: TDATA = 46'b0110101010000011111101100000000101011001011110;
        11'd845: TDATA = 46'b0110101001100011111001000000000011111110101010;
        11'd846: TDATA = 46'b0110101001000011110101000000000010100011111001;
        11'd847: TDATA = 46'b0110101000100011110100000000000001001001010011;
        11'd848: TDATA = 46'b0110101000000011110011111111111111011101100001;
        11'd849: TDATA = 46'b0110100111100011110100011111111100101000100110;
        11'd850: TDATA = 46'b0110100111000011110111011111111001110011111100;
        11'd851: TDATA = 46'b0110100110100011111010111111110110111111011001;
        11'd852: TDATA = 46'b0110100110000100000000011111110100001011000110;
        11'd853: TDATA = 46'b0110100101100100000110111111110001010110111100;
        11'd854: TDATA = 46'b0110100101000100001110111111101110100010111111;
        11'd855: TDATA = 46'b0110100100100100011000011111101011101111001110;
        11'd856: TDATA = 46'b0110100100000100100011011111101000111011101001;
        11'd857: TDATA = 46'b0110100011100100101111011111100110001000001111;
        11'd858: TDATA = 46'b0110100011000100111100111111100011010101000000;
        11'd859: TDATA = 46'b0110100010100101001011111111100000100001111110;
        11'd860: TDATA = 46'b0110100010000101011100011111011101101111001000;
        11'd861: TDATA = 46'b0110100001100101101101111111011010111100011100;
        11'd862: TDATA = 46'b0110100001000110000001011111011000001001111111;
        11'd863: TDATA = 46'b0110100000100110010101011111010101010111101001;
        11'd864: TDATA = 46'b0110100000000110101011111111010010100101100101;
        11'd865: TDATA = 46'b0110011111100111000011111111001111110011101101;
        11'd866: TDATA = 46'b0110011111000111011100011111001101000001111100;
        11'd867: TDATA = 46'b0110011110100111110110111111001010010000011010;
        11'd868: TDATA = 46'b0110011110001000010001111111000111011110111110;
        11'd869: TDATA = 46'b0110011101101000101101111111000100101101101101;
        11'd870: TDATA = 46'b0110011101001001001100111111000001111100110000;
        11'd871: TDATA = 46'b0110011100101001101100111110111111001011111100;
        11'd872: TDATA = 46'b0110011100001010001110111110111100011011011000;
        11'd873: TDATA = 46'b0110011011101010110000011110111001101010110100;
        11'd874: TDATA = 46'b0110011011001011010100011110110110111010100011;
        11'd875: TDATA = 46'b0110011010101011111001011110110100001010011011;
        11'd876: TDATA = 46'b0110011010001100100000011110110001011010100010;
        11'd877: TDATA = 46'b0110011001101101001000011110101110101010110010;
        11'd878: TDATA = 46'b0110011001001101110000111110101011111011001001;
        11'd879: TDATA = 46'b0110011000101110011100011110101001001011110101;
        11'd880: TDATA = 46'b0110011000001111001000011110100110011100100111;
        11'd881: TDATA = 46'b0110010111101111110101111110100011101101100110;
        11'd882: TDATA = 46'b0110010111010000100100111110100000111110110001;
        11'd883: TDATA = 46'b0110010110110001010100111110011110010000000101;
        11'd884: TDATA = 46'b0110010110010010000101111110011011100001100010;
        11'd885: TDATA = 46'b0110010101110010111000111110011000110011001111;
        11'd886: TDATA = 46'b0110010101010011101101011110010110000101001000;
        11'd887: TDATA = 46'b0110010100110100100011111110010011010111001111;
        11'd888: TDATA = 46'b0110010100010101011001111110010000101001011000;
        11'd889: TDATA = 46'b0110010011110110010010111110001101111011110101;
        11'd890: TDATA = 46'b0110010011010111001100111110001011001110011100;
        11'd891: TDATA = 46'b0110010010111000000111011110001000100001001001;
        11'd892: TDATA = 46'b0110010010011001000100011110000101110100001000;
        11'd893: TDATA = 46'b0110010001111010000000111110000011000111001000;
        11'd894: TDATA = 46'b0110010001011011000000011110000000011010011100;
        11'd895: TDATA = 46'b0110010000111100000000111101111101101101111010;
        11'd896: TDATA = 46'b0110010000011101000011011101111011000001100110;
        11'd897: TDATA = 46'b0110001111111110000101111101111000010101010111;
        11'd898: TDATA = 46'b0110001111011111001010111101110101101001011001;
        11'd899: TDATA = 46'b0110001111000000010000011101110010111101100001;
        11'd900: TDATA = 46'b0110001110100001010111011101110000010001110101;
        11'd901: TDATA = 46'b0110001110000010011111111101101101100110010110;
        11'd902: TDATA = 46'b0110001101100011101001011101101010111011000000;
        11'd903: TDATA = 46'b0110001101000100110100111101101000001111111000;
        11'd904: TDATA = 46'b0110001100100110000001111101100101100100111101;
        11'd905: TDATA = 46'b0110001100000111001111111101100010111010001011;
        11'd906: TDATA = 46'b0110001011101000011110111101100000001111100010;
        11'd907: TDATA = 46'b0110001011001001101111011101011101100101000101;
        11'd908: TDATA = 46'b0110001010101011000000111101011010111010110010;
        11'd909: TDATA = 46'b0110001010001100010100011101011000010000101101;
        11'd910: TDATA = 46'b0110001001101101101000011101010101100110101111;
        11'd911: TDATA = 46'b0110001001001110111111011101010010111101000101;
        11'd912: TDATA = 46'b0110001000110000010101111101010000010011011011;
        11'd913: TDATA = 46'b0110001000010001101110111101001101101010000100;
        11'd914: TDATA = 46'b0110000111110011001000011101001011000000110011;
        11'd915: TDATA = 46'b0110000111010100100011011101001000010111101101;
        11'd916: TDATA = 46'b0110000110110110000000011101000101101110110111;
        11'd917: TDATA = 46'b0110000110010111011101011101000011000110000100;
        11'd918: TDATA = 46'b0110000101111000111100111101000000011101100010;
        11'd919: TDATA = 46'b0110000101011010011100111100111101110101000111;
        11'd920: TDATA = 46'b0110000100111011111111011100111011001100111110;
        11'd921: TDATA = 46'b0110000100011101100010111100111000100100111101;
        11'd922: TDATA = 46'b0110000011111111000110111100110101111101000011;
        11'd923: TDATA = 46'b0110000011100000101011111100110011010101010010;
        11'd924: TDATA = 46'b0110000011000010010011011100110000101101110010;
        11'd925: TDATA = 46'b0110000010100011111011111100101110000110011100;
        11'd926: TDATA = 46'b0110000010000101100100111100101011011111001100;
        11'd927: TDATA = 46'b0110000001100111010000011100101000111000001101;
        11'd928: TDATA = 46'b0110000001001000111100011100100110010001010100;
        11'd929: TDATA = 46'b0110000000101010101001111100100011101010101000;
        11'd930: TDATA = 46'b0110000000001100011000011100100001000100000100;
        11'd931: TDATA = 46'b0101111111101110001000111100011110011101101111;
        11'd932: TDATA = 46'b0101111111001111111001111100011011110111100001;
        11'd933: TDATA = 46'b0101111110110001101100011100011001010001011110;
        11'd934: TDATA = 46'b0101111110010011100000011100010110101011100111;
        11'd935: TDATA = 46'b0101111101110101010101111100010100000101111100;
        11'd936: TDATA = 46'b0101111101010111001100111100010001100000011100;
        11'd937: TDATA = 46'b0101111100111001000100011100001110111011000011;
        11'd938: TDATA = 46'b0101111100011010111101011100001100010101110110;
        11'd939: TDATA = 46'b0101111011111100111000011100001001110000110111;
        11'd940: TDATA = 46'b0101111011011110110100011100000111001100000001;
        11'd941: TDATA = 46'b0101111011000000110000111100000100100111010010;
        11'd942: TDATA = 46'b0101111010100010101111111100000010000010110011;
        11'd943: TDATA = 46'b0101111010000100101111011011111111011110011011;
        11'd944: TDATA = 46'b0101111001100110110000011011111100111010001111;
        11'd945: TDATA = 46'b0101111001001000110010111011111010010110001111;
        11'd946: TDATA = 46'b0101111000101010110101011011110111110010010001;
        11'd947: TDATA = 46'b0101111000001100111001111011110101001110100011;
        11'd948: TDATA = 46'b0101110111101111000000011011110010101011000011;
        11'd949: TDATA = 46'b0101110111010001000111111011110000000111101011;
        11'd950: TDATA = 46'b0101110110110011001111111011101101100100011010;
        11'd951: TDATA = 46'b0101110110010101011001111011101011000001011000;
        11'd952: TDATA = 46'b0101110101110111100100111011101000011110011110;
        11'd953: TDATA = 46'b0101110101011001110001011011100101111011110000;
        11'd954: TDATA = 46'b0101110100111011111111011011100011011001001110;
        11'd955: TDATA = 46'b0101110100011110001101111011100000110110110001;
        11'd956: TDATA = 46'b0101110100000000011110111011011110010100100110;
        11'd957: TDATA = 46'b0101110011100010110000011011011011110010100001;
        11'd958: TDATA = 46'b0101110011000101000001111011011001010000100000;
        11'd959: TDATA = 46'b0101110010100111010111011011010110101110111000;
        11'd960: TDATA = 46'b0101110010001001101011111011010100001101001110;
        11'd961: TDATA = 46'b0101110001101100000010111011010001101011110100;
        11'd962: TDATA = 46'b0101110001001110011001111011001111001010011111;
        11'd963: TDATA = 46'b0101110000110000110011011011001100101001011010;
        11'd964: TDATA = 46'b0101110000010011001101011011001010001000011011;
        11'd965: TDATA = 46'b0101101111110101101000111011000111100111101000;
        11'd966: TDATA = 46'b0101101111011000000101011011000101000110111110;
        11'd967: TDATA = 46'b0101101110111010100100011011000010100110100101;
        11'd968: TDATA = 46'b0101101110011101000011111011000000000110010010;
        11'd969: TDATA = 46'b0101101101111111100011111010111101100110000101;
        11'd970: TDATA = 46'b0101101101100010000101111010111011000110000111;
        11'd971: TDATA = 46'b0101101101000100101000011010111000100110001110;
        11'd972: TDATA = 46'b0101101100100111001101011010110110000110100110;
        11'd973: TDATA = 46'b0101101100001001110010111010110011100111000101;
        11'd974: TDATA = 46'b0101101011101100011001011010110001000111101100;
        11'd975: TDATA = 46'b0101101011001111000000111010101110101000011100;
        11'd976: TDATA = 46'b0101101010110001101011011010101100001001100000;
        11'd977: TDATA = 46'b0101101010010100010101011010101001101010100101;
        11'd978: TDATA = 46'b0101101001110111000001011010100111001011110111;
        11'd979: TDATA = 46'b0101101001011001101110111010100100101101010101;
        11'd980: TDATA = 46'b0101101000111100011100111010100010001110111001;
        11'd981: TDATA = 46'b0101101000011111001011111010011111110000100110;
        11'd982: TDATA = 46'b0101101000000001111100111010011101010010100001;
        11'd983: TDATA = 46'b0101100111100100101101111010011010110100011111;
        11'd984: TDATA = 46'b0101100111000111100001011010011000010110101111;
        11'd985: TDATA = 46'b0101100110101010010101111010010101111001000111;
        11'd986: TDATA = 46'b0101100110001101001100011010010011011011101101;
        11'd987: TDATA = 46'b0101100101110000000011011010010000111110011001;
        11'd988: TDATA = 46'b0101100101010010111011011010001110100001001101;
        11'd989: TDATA = 46'b0101100100110101110100111010001100000100001110;
        11'd990: TDATA = 46'b0101100100011000101110111010001001100111010100;
        11'd991: TDATA = 46'b0101100011111011101010111010000111001010101000;
        11'd992: TDATA = 46'b0101100011011110101000011010000100101110001000;
        11'd993: TDATA = 46'b0101100011000001100101111010000010010001101011;
        11'd994: TDATA = 46'b0101100010100100100100111001111111110101011001;
        11'd995: TDATA = 46'b0101100010000111100101111001111101011001010101;
        11'd996: TDATA = 46'b0101100001101010101000011001111010111101011101;
        11'd997: TDATA = 46'b0101100001001101101011011001111000100001101011;
        11'd998: TDATA = 46'b0101100000110000101111011001110110000110000001;
        11'd999: TDATA = 46'b0101100000010011110101011001110011101010100110;
        11'd1000: TDATA = 46'b0101011111110110111100011001110001001111010011;
        11'd1001: TDATA = 46'b0101011111011010000011111001101110110100000110;
        11'd1002: TDATA = 46'b0101011110111101001100111001101100011001000100;
        11'd1003: TDATA = 46'b0101011110100000010111111001101001111110010000;
        11'd1004: TDATA = 46'b0101011110000011100011111001100111100011100101;
        11'd1005: TDATA = 46'b0101011101100110101111111001100101001000111101;
        11'd1006: TDATA = 46'b0101011101001001111101111001100010101110100011;
        11'd1007: TDATA = 46'b0101011100101101001101011001100000010100010101;
        11'd1008: TDATA = 46'b0101011100010000011101111001011101111010001111;
        11'd1009: TDATA = 46'b0101011011110011101111011001011011100000010001;
        11'd1010: TDATA = 46'b0101011011010111000001111001011001000110011100;
        11'd1011: TDATA = 46'b0101011010111010010101111001010110101100110011;
        11'd1012: TDATA = 46'b0101011010011101101011111001010100010011010111;
        11'd1013: TDATA = 46'b0101011010000001000001111001010001111001111111;
        11'd1014: TDATA = 46'b0101011001100100011001011001001111100000110001;
        11'd1015: TDATA = 46'b0101011001000111110010111001001101000111110010;
        11'd1016: TDATA = 46'b0101011000101011001100111001001010101110111000;
        11'd1017: TDATA = 46'b0101011000001110101000011001001000010110001010;
        11'd1018: TDATA = 46'b0101010111110010000100011001000101111101100010;
        11'd1019: TDATA = 46'b0101010111010101100001011001000011100101000010;
        11'd1020: TDATA = 46'b0101010110111001000000011001000001001100110000;
        11'd1021: TDATA = 46'b0101010110011100100000011000111110110100100110;
        11'd1022: TDATA = 46'b0101010110000000000010111000111100011100101101;
        11'd1023: TDATA = 46'b0101010101100011100100011000111010000100110010;
        11'd1024: TDATA = 46'b0101010101000111000111111000110111101101000101;
        11'd1025: TDATA = 46'b0101010100101010101100011000110101010101100000;
        11'd1026: TDATA = 46'b0101010100001110010010111000110010111110001001;
        11'd1027: TDATA = 46'b0101010011110001111001011000110000100110110101;
        11'd1028: TDATA = 46'b0101010011010101100001011000101110001111101100;
        11'd1029: TDATA = 46'b0101010010111001001011011000101011111000110001;
        11'd1030: TDATA = 46'b0101010010011100110101011000101001100001111010;
        11'd1031: TDATA = 46'b0101010010000000100001011000100111001011010000;
        11'd1032: TDATA = 46'b0101010001100100001110111000100100110100110001;
        11'd1033: TDATA = 46'b0101010001000111111100111000100010011110011000;
        11'd1034: TDATA = 46'b0101010000101011101100011000100000001000001001;
        11'd1035: TDATA = 46'b0101010000001111011100011000011101110010000001;
        11'd1036: TDATA = 46'b0101001111110011001101111000011011011100000100;
        11'd1037: TDATA = 46'b0101001111010111000001011000011001000110010101;
        11'd1038: TDATA = 46'b0101001110111010110101011000010110110000101011;
        11'd1039: TDATA = 46'b0101001110011110101010111000010100011011001100;
        11'd1040: TDATA = 46'b0101001110000010100000111000010010000101110011;
        11'd1041: TDATA = 46'b0101001101100110011000011000001111110000100110;
        11'd1042: TDATA = 46'b0101001101001010010001011000001101011011100011;
        11'd1043: TDATA = 46'b0101001100101110001010111000001011000110100110;
        11'd1044: TDATA = 46'b0101001100010010000101111000001000110001110100;
        11'd1045: TDATA = 46'b0101001011110110000001111000000110011101001010;
        11'd1046: TDATA = 46'b0101001011011001111111111000000100001000101110;
        11'd1047: TDATA = 46'b0101001010111101111101111000000001110100010101;
        11'd1048: TDATA = 46'b0101001010100001111101110111111111100000001010;
        11'd1049: TDATA = 46'b0101001010000101111110110111111101001100000111;
        11'd1050: TDATA = 46'b0101001001101010000000010111111010111000001010;
        11'd1051: TDATA = 46'b0101001001001110000011110111111000100100011010;
        11'd1052: TDATA = 46'b0101001000110010000111110111110110010000110001;
        11'd1053: TDATA = 46'b0101001000010110001101010111110011111101010010;
        11'd1054: TDATA = 46'b0101000111111010010100010111110001101001111110;
        11'd1055: TDATA = 46'b0101000111011110011011110111101111010110101111;
        11'd1056: TDATA = 46'b0101000111000010100100110111101101000011101100;
        11'd1057: TDATA = 46'b0101000110100110101111010111101010110000110100;
        11'd1058: TDATA = 46'b0101000110001010111001010111101000011101111100;
        11'd1059: TDATA = 46'b0101000101101111000110110111100110001011011001;
        11'd1060: TDATA = 46'b0101000101010011010011110111100011111000110111;
        11'd1061: TDATA = 46'b0101000100110111100001110111100001100110011101;
        11'd1062: TDATA = 46'b0101000100011011110001110111011111010100010001;
        11'd1063: TDATA = 46'b0101000100000000000010110111011101000010001101;
        11'd1064: TDATA = 46'b0101000011100100010100110111011010110000010001;
        11'd1065: TDATA = 46'b0101000011001000101000010111011000011110100001;
        11'd1066: TDATA = 46'b0101000010101100111100110111010110001100111000;
        11'd1067: TDATA = 46'b0101000010010001010001010111010011111011010010;
        11'd1068: TDATA = 46'b0101000001110101101000110111010001101010000000;
        11'd1069: TDATA = 46'b0101000001011010000000010111001111011000110000;
        11'd1070: TDATA = 46'b0101000000111110011001010111001101000111101011;
        11'd1071: TDATA = 46'b0101000000100010110011010111001010110110101110;
        11'd1072: TDATA = 46'b0101000000000111001101110111001000100101110111;
        11'd1073: TDATA = 46'b0100111111101011101010110111000110010101010000;
        11'd1074: TDATA = 46'b0100111111010000001000010111000100000100101110;
        11'd1075: TDATA = 46'b0100111110110100100110110111000001110100010101;
        11'd1076: TDATA = 46'b0100111110011001000101110110111111100100000010;
        11'd1077: TDATA = 46'b0100111101111101100111010110111101010011111110;
        11'd1078: TDATA = 46'b0100111101100010001000010110111011000011111011;
        11'd1079: TDATA = 46'b0100111101000110101011110110111000110100000111;
        11'd1080: TDATA = 46'b0100111100101011001111110110110110100100011010;
        11'd1081: TDATA = 46'b0100111100001111110101010110110100010100110111;
        11'd1082: TDATA = 46'b0100111011110100011011110110110010000101011100;
        11'd1083: TDATA = 46'b0100111011011001000011110110101111110110001100;
        11'd1084: TDATA = 46'b0100111010111101101011110110101101100110111111;
        11'd1085: TDATA = 46'b0100111010100010010101010110101011010111111101;
        11'd1086: TDATA = 46'b0100111010000111000000010110101001001001000110;
        11'd1087: TDATA = 46'b0100111001101011101100010110100110111010010110;
        11'd1088: TDATA = 46'b0100111001010000011001110110100100101011110010;
        11'd1089: TDATA = 46'b0100111000110101000111110110100010011101010011;
        11'd1090: TDATA = 46'b0100111000011001110111010110100000001110111110;
        11'd1091: TDATA = 46'b0100110111111110100111110110011110000000110010;
        11'd1092: TDATA = 46'b0100110111100011011000110110011011110010101011;
        11'd1093: TDATA = 46'b0100110111001000001011110110011001100100110010;
        11'd1094: TDATA = 46'b0100110110101100111111110110010111010111000001;
        11'd1095: TDATA = 46'b0100110110010001110100110110010101001001011000;
        11'd1096: TDATA = 46'b0100110101110110101010110110010010111011110111;
        11'd1097: TDATA = 46'b0100110101011011100001010110010000101110011011;
        11'd1098: TDATA = 46'b0100110101000000011001110110001110100001001101;
        11'd1099: TDATA = 46'b0100110100100101010011010110001100010100000111;
        11'd1100: TDATA = 46'b0100110100001010001101010110001010000111000110;
        11'd1101: TDATA = 46'b0100110011101111001000110110000111111010010000;
        11'd1102: TDATA = 46'b0100110011010100000101010110000101101101100010;
        11'd1103: TDATA = 46'b0100110010111001000011010110000011100000111110;
        11'd1104: TDATA = 46'b0100110010011110000001110110000001010100100001;
        11'd1105: TDATA = 46'b0100110010000011000001110101111111001000001101;
        11'd1106: TDATA = 46'b0100110001101000000010110101111100111100000010;
        11'd1107: TDATA = 46'b0100110001001101000100110101111010101111111111;
        11'd1108: TDATA = 46'b0100110000110010001000010101111000100100000110;
        11'd1109: TDATA = 46'b0100110000010111001100110101110110011000010110;
        11'd1110: TDATA = 46'b0100101111111100010001110101110100001100101011;
        11'd1111: TDATA = 46'b0100101111100001011000010101110010000001001010;
        11'd1112: TDATA = 46'b0100101111000110011111110101101111110101110010;
        11'd1113: TDATA = 46'b0100101110101011100111110101101101101010011111;
        11'd1114: TDATA = 46'b0100101110010000110001110101101011011111011001;
        11'd1115: TDATA = 46'b0100101101110101111100110101101001010100011011;
        11'd1116: TDATA = 46'b0100101101011011001000110101100111001001100101;
        11'd1117: TDATA = 46'b0100101101000000010101110101100100111110110111;
        11'd1118: TDATA = 46'b0100101100100101100011110101100010110100010001;
        11'd1119: TDATA = 46'b0100101100001010110010110101100000101001110011;
        11'd1120: TDATA = 46'b0100101011110000000011010101011110011111100000;
        11'd1121: TDATA = 46'b0100101011010101010100010101011100010101010010;
        11'd1122: TDATA = 46'b0100101010111010100110110101011010001011001111;
        11'd1123: TDATA = 46'b0100101010011111111001110101011000000001010000;
        11'd1124: TDATA = 46'b0100101010000101001111010101010101110111100010;
        11'd1125: TDATA = 46'b0100101001101010100100110101010011101101110110;
        11'd1126: TDATA = 46'b0100101001001111111011010101010001100100010011;
        11'd1127: TDATA = 46'b0100101000110101010010110101001111011010110111;
        11'd1128: TDATA = 46'b0100101000011010101011110101001101010001100110;
        11'd1129: TDATA = 46'b0100101000000000000101010101001011001000011010;
        11'd1130: TDATA = 46'b0100100111100101100000110101001000111111011011;
        11'd1131: TDATA = 46'b0100100111001010111100010101000110110110011111;
        11'd1132: TDATA = 46'b0100100110110000011001010101000100101101101101;
        11'd1133: TDATA = 46'b0100100110010101111000010101000010100101001001;
        11'd1134: TDATA = 46'b0100100101111011010110110101000000011100100100;
        11'd1135: TDATA = 46'b0100100101100000110111110100111110010100010000;
        11'd1136: TDATA = 46'b0100100101000110011000010100111100001011111011;
        11'd1137: TDATA = 46'b0100100100101011111011010100111010000011110110;
        11'd1138: TDATA = 46'b0100100100010001011110110100110111111011110110;
        11'd1139: TDATA = 46'b0100100011110111000011010100110101110011111111;
        11'd1140: TDATA = 46'b0100100011011100101000110100110011101100001111;
        11'd1141: TDATA = 46'b0100100011000010001111010100110001100100100111;
        11'd1142: TDATA = 46'b0100100010100111110111010100101111011101001001;
        11'd1143: TDATA = 46'b0100100010001101011111110100101101010101110001;
        11'd1144: TDATA = 46'b0100100001110011001001110100101011001110100011;
        11'd1145: TDATA = 46'b0100100001011000110100110100101001000111011100;
        11'd1146: TDATA = 46'b0100100000111110100000110100100111000000011110;
        11'd1147: TDATA = 46'b0100100000100100001101110100100100111001101000;
        11'd1148: TDATA = 46'b0100100000001001111100010100100010110010111100;
        11'd1149: TDATA = 46'b0100011111101111101011010100100000101100010101;
        11'd1150: TDATA = 46'b0100011111010101011011010100011110100101110110;
        11'd1151: TDATA = 46'b0100011110111011001100010100011100011111011111;
        11'd1152: TDATA = 46'b0100011110100000111110110100011010011001010010;
        11'd1153: TDATA = 46'b0100011110000110110001110100011000010011001010;
        11'd1154: TDATA = 46'b0100011101101100100110110100010110001101010000;
        11'd1155: TDATA = 46'b0100011101010010011011110100010100000111011000;
        11'd1156: TDATA = 46'b0100011100111000010010110100010010000001101101;
        11'd1157: TDATA = 46'b0100011100011110001001110100001111111100000100;
        11'd1158: TDATA = 46'b0100011100000100000001110100001101110110100100;
        11'd1159: TDATA = 46'b0100011011101001111100010100001011110001010011;
        11'd1160: TDATA = 46'b0100011011001111110110110100001001101100000100;
        11'd1161: TDATA = 46'b0100011010110101110001110100000111100110111011;
        11'd1162: TDATA = 46'b0100011010011011101111010100000101100010000001;
        11'd1163: TDATA = 46'b0100011010000001101100110100000011011101001010;
        11'd1164: TDATA = 46'b0100011001100111101011110100000001011000011101;
        11'd1165: TDATA = 46'b0100011001001101101011110011111111010011110111;
        11'd1166: TDATA = 46'b0100011000110011101100010011111101001111010111;
        11'd1167: TDATA = 46'b0100011000011001101101110011111011001010111111;
        11'd1168: TDATA = 46'b0100010111111111110000110011111001000110110001;
        11'd1169: TDATA = 46'b0100010111100101110100110011110111000010101011;
        11'd1170: TDATA = 46'b0100010111001011111001110011110100111110101100;
        11'd1171: TDATA = 46'b0100010110110010000000010011110010111010111000;
        11'd1172: TDATA = 46'b0100010110011000000111010011110000110111001001;
        11'd1173: TDATA = 46'b0100010101111110001111010011101110110011100001;
        11'd1174: TDATA = 46'b0100010101100100010111110011101100101111111111;
        11'd1175: TDATA = 46'b0100010101001010100010110011101010101100101100;
        11'd1176: TDATA = 46'b0100010100110000101101010011101000101001011001;
        11'd1177: TDATA = 46'b0100010100010110111001110011100110100110010011;
        11'd1178: TDATA = 46'b0100010011111101000111010011100100100011010101;
        11'd1179: TDATA = 46'b0100010011100011010100110011100010100000011001;
        11'd1180: TDATA = 46'b0100010011001001100100010011100000011101101010;
        11'd1181: TDATA = 46'b0100010010101111110100010011011110011011000000;
        11'd1182: TDATA = 46'b0100010010010110000101110011011100011000100000;
        11'd1183: TDATA = 46'b0100010001111100011000010011011010010110001000;
        11'd1184: TDATA = 46'b0100010001100010101011110011011000010011110111;
        11'd1185: TDATA = 46'b0100010001001000111111110011010110010001101100;
        11'd1186: TDATA = 46'b0100010000101111010101010011010100001111101011;
        11'd1187: TDATA = 46'b0100010000010101101011110011010010001101110001;
        11'd1188: TDATA = 46'b0100001111111100000011010011010000001011111111;
        11'd1189: TDATA = 46'b0100001111100010011011110011001110001010010101;
        11'd1190: TDATA = 46'b0100001111001000110101010011001100001000110010;
        11'd1191: TDATA = 46'b0100001110101111001111010011001010000111010101;
        11'd1192: TDATA = 46'b0100001110010101101011010011001000000110000100;
        11'd1193: TDATA = 46'b0100001101111100000111010011000110000100110101;
        11'd1194: TDATA = 46'b0100001101100010100100110011000100000011110001;
        11'd1195: TDATA = 46'b0100001101001001000011110011000010000010110111;
        11'd1196: TDATA = 46'b0100001100101111100010110011000000000010000000;
        11'd1197: TDATA = 46'b0100001100010110000011110010111110000001010101;
        11'd1198: TDATA = 46'b0100001011111100100100010010111100000000101010;
        11'd1199: TDATA = 46'b0100001011100011000111010010111010000000001110;
        11'd1200: TDATA = 46'b0100001011001001101010110010110111111111110111;
        11'd1201: TDATA = 46'b0100001010110000001111010010110101111111101000;
        11'd1202: TDATA = 46'b0100001010010110110100110010110011111111100001;
        11'd1203: TDATA = 46'b0100001001111101011011010010110001111111100001;
        11'd1204: TDATA = 46'b0100001001100100000010110010101111111111101000;
        11'd1205: TDATA = 46'b0100001001001010101011010010101101111111110111;
        11'd1206: TDATA = 46'b0100001000110001010100110010101100000000001110;
        11'd1207: TDATA = 46'b0100001000010111111111010010101010000000101100;
        11'd1208: TDATA = 46'b0100000111111110101011010010101000000001010100;
        11'd1209: TDATA = 46'b0100000111100101010111010010100110000001111111;
        11'd1210: TDATA = 46'b0100000111001100000100110010100100000010110100;
        11'd1211: TDATA = 46'b0100000110110010110011010010100010000011110000;
        11'd1212: TDATA = 46'b0100000110011001100010110010100000000100110100;
        11'd1213: TDATA = 46'b0100000110000000010011010010011110000101111111;
        11'd1214: TDATA = 46'b0100000101100111000100110010011100000111010010;
        11'd1215: TDATA = 46'b0100000101001101110111010010011010001000101101;
        11'd1216: TDATA = 46'b0100000100110100101001110010011000001010001010;
        11'd1217: TDATA = 46'b0100000100011011011111010010010110001011111000;
        11'd1218: TDATA = 46'b0100000100000010010100010010010100001101100110;
        11'd1219: TDATA = 46'b0100000011101001001010110010010010001111011111;
        11'd1220: TDATA = 46'b0100000011010000000001110010010000010001011100;
        11'd1221: TDATA = 46'b0100000010110110111010110010001110010011100110;
        11'd1222: TDATA = 46'b0100000010011101110011110010001100010101110010;
        11'd1223: TDATA = 46'b0100000010000100101101110010001010011000000110;
        11'd1224: TDATA = 46'b0100000001101011101001010010001000011010100100;
        11'd1225: TDATA = 46'b0100000001010010100101010010000110011101000110;
        11'd1226: TDATA = 46'b0100000000111001100010110010000100011111110011;
        11'd1227: TDATA = 46'b0100000000100000100000110010000010100010100101;
        11'd1228: TDATA = 46'b0100000000000111100000010010000000100101100000;
        11'd1229: TDATA = 46'b0011111111101110100000010001111110101000100001;
        11'd1230: TDATA = 46'b0011111111010101100001010001111100101011101001;
        11'd1231: TDATA = 46'b0011111110111100100011110001111010101110111010;
        11'd1232: TDATA = 46'b0011111110100011100111010001111000110010010100;
        11'd1233: TDATA = 46'b0011111110001010101011010001110110110101110010;
        11'd1234: TDATA = 46'b0011111101110001110000010001110100111001011000;
        11'd1235: TDATA = 46'b0011111101011000110110110001110010111101000111;
        11'd1236: TDATA = 46'b0011111100111111111101010001110001000000111001;
        11'd1237: TDATA = 46'b0011111100100111000101010001101111000100110101;
        11'd1238: TDATA = 46'b0011111100001110001101110001101101001000110110;
        11'd1239: TDATA = 46'b0011111011110101010111110001101011001101000000;
        11'd1240: TDATA = 46'b0011111011011100100011010001101001010001010101;
        11'd1241: TDATA = 46'b0011111011000011101111010001100111010101101110;
        11'd1242: TDATA = 46'b0011111010101010111011110001100101011010001101;
        11'd1243: TDATA = 46'b0011111010010010001001110001100011011110110101;
        11'd1244: TDATA = 46'b0011111001111001011000010001100001100011100010;
        11'd1245: TDATA = 46'b0011111001100000100111110001011111101000010110;
        11'd1246: TDATA = 46'b0011111001000111111000010001011101101101010010;
        11'd1247: TDATA = 46'b0011111000101111001001110001011011110010010110;
        11'd1248: TDATA = 46'b0011111000010110011100110001011001110111100011;
        11'd1249: TDATA = 46'b0011110111111101110000010001010111111100110101;
        11'd1250: TDATA = 46'b0011110111100101000100110001010110000010001110;
        11'd1251: TDATA = 46'b0011110111001100011010110001010100000111110001;
        11'd1252: TDATA = 46'b0011110110110011110000110001010010001101010110;
        11'd1253: TDATA = 46'b0011110110011011000111110001010000010011000011;
        11'd1254: TDATA = 46'b0011110110000010100000010001001110011000111010;
        11'd1255: TDATA = 46'b0011110101101001111001010001001100011110110101;
        11'd1256: TDATA = 46'b0011110101010001010011110001001010100100111010;
        11'd1257: TDATA = 46'b0011110100111000101111010001001000101011000111;
        11'd1258: TDATA = 46'b0011110100100000001011010001000110110001011001;
        11'd1259: TDATA = 46'b0011110100000111101000010001000100110111110001;
        11'd1260: TDATA = 46'b0011110011101111000101110001000010111110001111;
        11'd1261: TDATA = 46'b0011110011010110100100110001000001000100110110;
        11'd1262: TDATA = 46'b0011110010111110000100110000111111001011100101;
        11'd1263: TDATA = 46'b0011110010100101100101110000111101010010011011;
        11'd1264: TDATA = 46'b0011110010001101001000010000111011011001011010;
        11'd1265: TDATA = 46'b0011110001110100101010110000111001100000011100;
        11'd1266: TDATA = 46'b0011110001011100001110110000110111100111101000;
        11'd1267: TDATA = 46'b0011110001000011110011010000110101101110111001;
        11'd1268: TDATA = 46'b0011110000101011011000010000110011110110001110;
        11'd1269: TDATA = 46'b0011110000010010111111010000110001111101110000;
        11'd1270: TDATA = 46'b0011101111111010100110110000110000000101010110;
        11'd1271: TDATA = 46'b0011101111100010001111010000101110001101000100;
        11'd1272: TDATA = 46'b0011101111001001111000010000101100010100110110;
        11'd1273: TDATA = 46'b0011101110110001100011010000101010011100110101;
        11'd1274: TDATA = 46'b0011101110011001001101110000101000100100110011;
        11'd1275: TDATA = 46'b0011101110000000111010110000100110101101000000;
        11'd1276: TDATA = 46'b0011101101101000100111010000100100110101001101;
        11'd1277: TDATA = 46'b0011101101010000010101010000100010111101100100;
        11'd1278: TDATA = 46'b0011101100111000000100010000100001000110000010;
        11'd1279: TDATA = 46'b0011101100011111110100010000011111001110100111;
        11'd1280: TDATA = 46'b0011101100000111100101010000011101010111010011;
        11'd1281: TDATA = 46'b0011101011101111010110110000011011100000000100;
        11'd1282: TDATA = 46'b0011101011010111001001010000011001101000111101;
        11'd1283: TDATA = 46'b0011101010111110111101010000010111110001111110;
        11'd1284: TDATA = 46'b0011101010100110110001010000010101111011000011;
        11'd1285: TDATA = 46'b0011101010001110100111010000010100000100010011;
        11'd1286: TDATA = 46'b0011101001110110011101110000010010001101101000;
        11'd1287: TDATA = 46'b0011101001011110010100110000010000010111000010;
        11'd1288: TDATA = 46'b0011101001000110001101010000001110100000100101;
        11'd1289: TDATA = 46'b0011101000101110000110110000001100101010010000;
        11'd1290: TDATA = 46'b0011101000010110000000110000001010110011111111;
        11'd1291: TDATA = 46'b0011100111111101111011110000001000111101110110;
        11'd1292: TDATA = 46'b0011100111100101110111110000000111000111110100;
        11'd1293: TDATA = 46'b0011100111001101110100010000000101010001110110;
        11'd1294: TDATA = 46'b0011100110110101110010110000000011011100000101;
        11'd1295: TDATA = 46'b0011100110011101110000110000000001100110010011;
        11'd1296: TDATA = 46'b0011100110000101110000101111111111110000101101;
        11'd1297: TDATA = 46'b0011100101101101110001001111111101111011001100;
        11'd1298: TDATA = 46'b0011100101010101110011001111111100000101110101;
        11'd1299: TDATA = 46'b0011100100111101110101001111111010010000100000;
        11'd1300: TDATA = 46'b0011100100100101111000101111111000011011010100;
        11'd1301: TDATA = 46'b0011100100001101111100101111110110100110001101;
        11'd1302: TDATA = 46'b0011100011110110000010101111110100110001010010;
        11'd1303: TDATA = 46'b0011100011011110001000001111110010111100010111;
        11'd1304: TDATA = 46'b0011100011000110001111001111110001000111100110;
        11'd1305: TDATA = 46'b0011100010101110010111001111101111010010111100;
        11'd1306: TDATA = 46'b0011100010010110011111101111101101011110010110;
        11'd1307: TDATA = 46'b0011100001111110101001001111101011101001110111;
        11'd1308: TDATA = 46'b0011100001100110110100001111101001110101100010;
        11'd1309: TDATA = 46'b0011100001001111000000001111101000000001010100;
        11'd1310: TDATA = 46'b0011100000110111001100001111100110001101001000;
        11'd1311: TDATA = 46'b0011100000011111011001101111100100011001000110;
        11'd1312: TDATA = 46'b0011100000000111101000001111100010100101001011;
        11'd1313: TDATA = 46'b0011011111101111110111001111100000110001010101;
        11'd1314: TDATA = 46'b0011011111011000000111001111011110111101100101;
        11'd1315: TDATA = 46'b0011011111000000011000001111011101001001111101;
        11'd1316: TDATA = 46'b0011011110101000101001101111011011010110011001;
        11'd1317: TDATA = 46'b0011011110010000111100001111011001100010111101;
        11'd1318: TDATA = 46'b0011011101111001010000001111010111101111101001;
        11'd1319: TDATA = 46'b0011011101100001100100101111010101111100011011;
        11'd1320: TDATA = 46'b0011011101001001111010101111010100001001010110;
        11'd1321: TDATA = 46'b0011011100110010010000101111010010010110010011;
        11'd1322: TDATA = 46'b0011011100011010101000001111010000100011011010;
        11'd1323: TDATA = 46'b0011011100000011000000001111001110110000100101;
        11'd1324: TDATA = 46'b0011011011101011011001001111001100111101110111;
        11'd1325: TDATA = 46'b0011011011010011110011001111001011001011010001;
        11'd1326: TDATA = 46'b0011011010111100001101101111001001011000101111;
        11'd1327: TDATA = 46'b0011011010100100101001101111000111100110010110;
        11'd1328: TDATA = 46'b0011011010001101000110101111000101110100000100;
        11'd1329: TDATA = 46'b0011011001110101100100001111000100000001110111;
        11'd1330: TDATA = 46'b0011011001011110000010101111000010001111110001;
        11'd1331: TDATA = 46'b0011011001000110100001101111000000011101110000;
        11'd1332: TDATA = 46'b0011011000101111000001101110111110101011110110;
        11'd1333: TDATA = 46'b0011011000010111100011101110111100111010000111;
        11'd1334: TDATA = 46'b0011011000000000000100101110111011001000010110;
        11'd1335: TDATA = 46'b0011010111101000101000001110111001010110110011;
        11'd1336: TDATA = 46'b0011010111010001001011101110110111100101010010;
        11'd1337: TDATA = 46'b0011010110111001110000101110110101110011111011;
        11'd1338: TDATA = 46'b0011010110100010010101101110110100000010100101;
        11'd1339: TDATA = 46'b0011010110001010111100001110110010010001011001;
        11'd1340: TDATA = 46'b0011010101110011100011101110110000100000010100;
        11'd1341: TDATA = 46'b0011010101011100001011101110101110101111010100;
        11'd1342: TDATA = 46'b0011010101000100110100101110101100111110011011;
        11'd1343: TDATA = 46'b0011010100101101011111001110101011001101101011;
        11'd1344: TDATA = 46'b0011010100010110001001001110101001011100111010;
        11'd1345: TDATA = 46'b0011010011111110110101001110100111101100010110;
        11'd1346: TDATA = 46'b0011010011100111100010101110100101111011111011;
        11'd1347: TDATA = 46'b0011010011010000001111101110100100001011011111;
        11'd1348: TDATA = 46'b0011010010111000111101101110100010011011001011;
        11'd1349: TDATA = 46'b0011010010100001101101001110100000101011000000;
        11'd1350: TDATA = 46'b0011010010001010011101001110011110111010111001;
        11'd1351: TDATA = 46'b0011010001110011001101101110011101001010110111;
        11'd1352: TDATA = 46'b0011010001011100000000001110011011011011000001;
        11'd1353: TDATA = 46'b0011010001000100110010101110011001101011001100;
        11'd1354: TDATA = 46'b0011010000101101100101101110010111111011011101;
        11'd1355: TDATA = 46'b0011010000010110011011001110010110001011111011;
        11'd1356: TDATA = 46'b0011001111111111010000001110010100011100011001;
        11'd1357: TDATA = 46'b0011001111101000000110101110010010101101000000;
        11'd1358: TDATA = 46'b0011001111010000111101101110010000111101101100;
        11'd1359: TDATA = 46'b0011001110111001110101001110001111001110011101;
        11'd1360: TDATA = 46'b0011001110100010101101101110001101011111010100;
        11'd1361: TDATA = 46'b0011001110001011101000001110001011110000010111;
        11'd1362: TDATA = 46'b0011001101110100100010101110001010000001011100;
        11'd1363: TDATA = 46'b0011001101011101011101101110001000010010100110;
        11'd1364: TDATA = 46'b0011001101000110011001101110000110100011110110;
        11'd1365: TDATA = 46'b0011001100101111010111101110000100110101010010;
        11'd1366: TDATA = 46'b0011001100011000010100101110000011000110101011;
        11'd1367: TDATA = 46'b0011001100000001010100001110000001011000010011;
        11'd1368: TDATA = 46'b0011001011101010010011101101111111101001111100;
        11'd1369: TDATA = 46'b0011001011010011010100001101111101111011101101;
        11'd1370: TDATA = 46'b0011001010111100010101101101111100001101100100;
        11'd1371: TDATA = 46'b0011001010100101011000001101111010011111100010;
        11'd1372: TDATA = 46'b0011001010001110011011101101111000110001100111;
        11'd1373: TDATA = 46'b0011001001110111011111101101110111000011110000;
        11'd1374: TDATA = 46'b0011001001100000100100101101110101010110000001;
        11'd1375: TDATA = 46'b0011001001001001101010101101110011101000011000;
        11'd1376: TDATA = 46'b0011001000110010110000101101110001111010110001;
        11'd1377: TDATA = 46'b0011001000011011111000001101110000001101010011;
        11'd1378: TDATA = 46'b0011001000000101000000001101101110011111111010;
        11'd1379: TDATA = 46'b0011000111101110001001101101101100110010101010;
        11'd1380: TDATA = 46'b0011000111010111010011101101101011000101011110;
        11'd1381: TDATA = 46'b0011000111000000011111001101101001011000011100;
        11'd1382: TDATA = 46'b0011000110101001101010101101100111101011011100;
        11'd1383: TDATA = 46'b0011000110010010110111001101100101111110100010;
        11'd1384: TDATA = 46'b0011000101111100000100001101100100010001101101;
        11'd1385: TDATA = 46'b0011000101100101010010101101100010100101000001;
        11'd1386: TDATA = 46'b0011000101001110100001101101100000111000011010;
        11'd1387: TDATA = 46'b0011000100110111110001101101011111001011111001;
        11'd1388: TDATA = 46'b0011000100100001000010101101011101011111011111;
        11'd1389: TDATA = 46'b0011000100001010010100001101011011110011001010;
        11'd1390: TDATA = 46'b0011000011110011100111001101011010000110111101;
        11'd1391: TDATA = 46'b0011000011011100111001101101011000011010110000;
        11'd1392: TDATA = 46'b0011000011000110001111001101010110101110110100;
        11'd1393: TDATA = 46'b0011000010101111100011101101010101000010110101;
        11'd1394: TDATA = 46'b0011000010011000111001001101010011010110111100;
        11'd1395: TDATA = 46'b0011000010000010010000101101010001101011010000;
        11'd1396: TDATA = 46'b0011000001101011100111101101001111111111100010;
        11'd1397: TDATA = 46'b0011000001010101000000001101001110010011111110;
        11'd1398: TDATA = 46'b0011000000111110011001001101001100101000011110;
        11'd1399: TDATA = 46'b0011000000100111110011101101001010111101001000;
        11'd1400: TDATA = 46'b0011000000010001001110101101001001010001110101;
        11'd1401: TDATA = 46'b0010111111111010101001101101000111100110100101;
        11'd1402: TDATA = 46'b0010111111100100000111001101000101111011100011;
        11'd1403: TDATA = 46'b0010111111001101100100001101000100010000100000;
        11'd1404: TDATA = 46'b0010111110110111000010101101000010100101100110;
        11'd1405: TDATA = 46'b0010111110100000100001101101000000111010110001;
        11'd1406: TDATA = 46'b0010111110001010000001101100111111010000000010;
        11'd1407: TDATA = 46'b0010111101110011100010101100111101100101011010;
        11'd1408: TDATA = 46'b0010111101011101000100001100111011111010110111;
        11'd1409: TDATA = 46'b0010111101000110100110101100111010010000011010;
        11'd1410: TDATA = 46'b0010111100110000001001101100111000100110000010;
        11'd1411: TDATA = 46'b0010111100011001101101101100110110111011110000;
        11'd1412: TDATA = 46'b0010111100000011010011001100110101010001100111;
        11'd1413: TDATA = 46'b0010111011101100111000001100110011100111011110;
        11'd1414: TDATA = 46'b0010111011010110011111001100110001111101100000;
        11'd1415: TDATA = 46'b0010111011000000000110101100110000010011100111;
        11'd1416: TDATA = 46'b0010111010101001101111001100101110101001110100;
        11'd1417: TDATA = 46'b0010111010010011010111101100101101000000000011;
        11'd1418: TDATA = 46'b0010111001111101000001101100101011010110011100;
        11'd1419: TDATA = 46'b0010111001100110101100101100101001101100111011;
        11'd1420: TDATA = 46'b0010111001010000011000001100101000000011011110;
        11'd1421: TDATA = 46'b0010111000111010000100101100100110011010001000;
        11'd1422: TDATA = 46'b0010111000100011110001101100100100110000110110;
        11'd1423: TDATA = 46'b0010111000001101100000001100100011000111101101;
        11'd1424: TDATA = 46'b0010110111110111001110101100100001011110100111;
        11'd1425: TDATA = 46'b0010110111100000111110101100011111110101101001;
        11'd1426: TDATA = 46'b0010110111001010101111001100011110001100101111;
        11'd1427: TDATA = 46'b0010110110110100100000001100011100100011111010;
        11'd1428: TDATA = 46'b0010110110011110010001101100011010111011001001;
        11'd1429: TDATA = 46'b0010110110001000000101001100011001010010100100;
        11'd1430: TDATA = 46'b0010110101110001111001001100010111101010000010;
        11'd1431: TDATA = 46'b0010110101011011101101001100010110000001100011;
        11'd1432: TDATA = 46'b0010110101000101100011001100010100011001001111;
        11'd1433: TDATA = 46'b0010110100101111011001001100010010110000111101;
        11'd1434: TDATA = 46'b0010110100011001010000101100010001001000110100;
        11'd1435: TDATA = 46'b0010110100000011001000001100001111100000101101;
        11'd1436: TDATA = 46'b0010110011101101000001001100001101111000101110;
        11'd1437: TDATA = 46'b0010110011010110111001101100001100010000110000;
        11'd1438: TDATA = 46'b0010110011000000110100101100001010101000111111;
        11'd1439: TDATA = 46'b0010110010101010101111101100001001000001010000;
        11'd1440: TDATA = 46'b0010110010010100101011101100000111011001100111;
        11'd1441: TDATA = 46'b0010110001111110101000001100000101110010000011;
        11'd1442: TDATA = 46'b0010110001101000100101001100000100001010100011;
        11'd1443: TDATA = 46'b0010110001010010100100001100000010100011001110;
        11'd1444: TDATA = 46'b0010110000111100100011101100000000111011111110;
        11'd1445: TDATA = 46'b0010110000100110100011101011111111010100110001;
        11'd1446: TDATA = 46'b0010110000010000100011101011111101101101100111;
        11'd1447: TDATA = 46'b0010101111111010100101101011111100000110101000;
        11'd1448: TDATA = 46'b0010101111100100100111101011111010011111101011;
        11'd1449: TDATA = 46'b0010101111001110101011001011111000111000110110;
        11'd1450: TDATA = 46'b0010101110111000101110101011110111010010000100;
        11'd1451: TDATA = 46'b0010101110100010110011101011110101101011011010;
        11'd1452: TDATA = 46'b0010101110001100111001001011110100000100110101;
        11'd1453: TDATA = 46'b0010101101110110111111001011110010011110010100;
        11'd1454: TDATA = 46'b0010101101100001000110101011110000110111111100;
        11'd1455: TDATA = 46'b0010101101001011001110101011101111010001101000;
        11'd1456: TDATA = 46'b0010101100110101010111101011101101101011011010;
        11'd1457: TDATA = 46'b0010101100011111100001001011101100000101010001;
        11'd1458: TDATA = 46'b0010101100001001101011001011101010011111001100;
        11'd1459: TDATA = 46'b0010101011110011110111001011101000111001010010;
        11'd1460: TDATA = 46'b0010101011011110000010101011100111010011011000;
        11'd1461: TDATA = 46'b0010101011001000001111001011100101101101100100;
        11'd1462: TDATA = 46'b0010101010110010011100101011100100000111110111;
        11'd1463: TDATA = 46'b0010101010011100101011001011100010100010010000;
        11'd1464: TDATA = 46'b0010101010000110111010101011100000111100110000;
        11'd1465: TDATA = 46'b0010101001110001001010101011011111010111010100;
        11'd1466: TDATA = 46'b0010101001011011011010101011011101110001111010;
        11'd1467: TDATA = 46'b0010101001000101101100001011011100001100101000;
        11'd1468: TDATA = 46'b0010101000101111111110101011011010100111011110;
        11'd1469: TDATA = 46'b0010101000011010010001001011011001000010010101;
        11'd1470: TDATA = 46'b0010101000000100100101001011010111011101010100;
        11'd1471: TDATA = 46'b0010100111101110111010101011010101111000011101;
        11'd1472: TDATA = 46'b0010100111011001001111101011010100010011100101;
        11'd1473: TDATA = 46'b0010100111000011100101101011010010101110110100;
        11'd1474: TDATA = 46'b0010100110101101111100101011010001001010001001;
        11'd1475: TDATA = 46'b0010100110011000010100101011001111100101100100;
        11'd1476: TDATA = 46'b0010100110000010101101001011001110000001000100;
        11'd1477: TDATA = 46'b0010100101101101000110101011001100011100101010;
        11'd1478: TDATA = 46'b0010100101010111100000101011001010111000010101;
        11'd1479: TDATA = 46'b0010100101000001111011101011001001010100000110;
        11'd1480: TDATA = 46'b0010100100101100010111101011000111101111111101;
        11'd1481: TDATA = 46'b0010100100010110110100001011000110001011111000;
        11'd1482: TDATA = 46'b0010100100000001010001001011000100100111111000;
        11'd1483: TDATA = 46'b0010100011101011110000001011000011000100000011;
        11'd1484: TDATA = 46'b0010100011010110001101101011000001100000001000;
        11'd1485: TDATA = 46'b0010100011000000101101101010111111111100011011;
        11'd1486: TDATA = 46'b0010100010101011001110101010111110011000110100;
        11'd1487: TDATA = 46'b0010100010010101101111101010111100110101001111;
        11'd1488: TDATA = 46'b0010100010000000010001101010111011010001110001;
        11'd1489: TDATA = 46'b0010100001101010110100001010111001101110010111;
        11'd1490: TDATA = 46'b0010100001010101010111101010111000001011000011;
        11'd1491: TDATA = 46'b0010100000111111111011101010110110100111110011;
        11'd1492: TDATA = 46'b0010100000101010100001001010110101000100101100;
        11'd1493: TDATA = 46'b0010100000010101000111001010110011100001101001;
        11'd1494: TDATA = 46'b0010011111111111101101101010110001111110101010;
        11'd1495: TDATA = 46'b0010011111101010010101001010110000011011110010;
        11'd1496: TDATA = 46'b0010011111010100111101001010101110111000111110;
        11'd1497: TDATA = 46'b0010011110111111100101101010101101010110001110;
        11'd1498: TDATA = 46'b0010011110101010001111101010101011110011100110;
        11'd1499: TDATA = 46'b0010011110010100111010101010101010010001000101;
        11'd1500: TDATA = 46'b0010011101111111100101101010101000101110100110;
        11'd1501: TDATA = 46'b0010011101101010010001001010100111001100001010;
        11'd1502: TDATA = 46'b0010011101010100111110101010100101101001111010;
        11'd1503: TDATA = 46'b0010011100111111101100001010100100000111101100;
        11'd1504: TDATA = 46'b0010011100101010011010101010100010100101100100;
        11'd1505: TDATA = 46'b0010011100010101001001001010100001000011011101;
        11'd1506: TDATA = 46'b0010011011111111111001001010011111100001100000;
        11'd1507: TDATA = 46'b0010011011101010101001101010011101111111100110;
        11'd1508: TDATA = 46'b0010011011010101011011101010011100011101110101;
        11'd1509: TDATA = 46'b0010011011000000001101101010011010111100000110;
        11'd1510: TDATA = 46'b0010011010101011000000001010011001011010011011;
        11'd1511: TDATA = 46'b0010011010010101110100001010010111111000111001;
        11'd1512: TDATA = 46'b0010011010000000101000001010010110010111011000;
        11'd1513: TDATA = 46'b0010011001101011011101001010010100110101111110;
        11'd1514: TDATA = 46'b0010011001010110010011101010010011010100101100;
        11'd1515: TDATA = 46'b0010011001000001001010101010010001110011011111;
        11'd1516: TDATA = 46'b0010011000101100000001101010010000010010010011;
        11'd1517: TDATA = 46'b0010011000010110111001101010001110110001001101;
        11'd1518: TDATA = 46'b0010011000000001110011001010001101010000010000;
        11'd1519: TDATA = 46'b0010010111101100101100101010001011101111010101;
        11'd1520: TDATA = 46'b0010010111010111100111001010001010001110100000;
        11'd1521: TDATA = 46'b0010010111000010100011001010001000101101110100;
        11'd1522: TDATA = 46'b0010010110101101011111001010000111001101001010;
        11'd1523: TDATA = 46'b0010010110011000011011101010000101101100100011;
        11'd1524: TDATA = 46'b0010010110000011011000101010000100001100000001;
        11'd1525: TDATA = 46'b0010010101101110010111001010000010101011100111;
        11'd1526: TDATA = 46'b0010010101011001010101101010000001001011001111;
        11'd1527: TDATA = 46'b0010010101000100010101101001111111101011000000;
        11'd1528: TDATA = 46'b0010010100101111010110101001111110001010110110;
        11'd1529: TDATA = 46'b0010010100011010011000001001111100101010110001;
        11'd1530: TDATA = 46'b0010010100000101011001101001111011001010101110;
        11'd1531: TDATA = 46'b0010010011110000011100101001111001101010110011;
        11'd1532: TDATA = 46'b0010010011011011100000001001111000001010111100;
        11'd1533: TDATA = 46'b0010010011000110100100101001110110101011001100;
        11'd1534: TDATA = 46'b0010010010110001101001001001110101001011011101;
        11'd1535: TDATA = 46'b0010010010011100101111001001110011101011110110;
        11'd1536: TDATA = 46'b0010010010000111110101101001110010001100010100;
        11'd1537: TDATA = 46'b0010010001110010111101001001110000101100111000;
        11'd1538: TDATA = 46'b0010010001011110000101001001101111001101100000;
        11'd1539: TDATA = 46'b0010010001001001001101101001101101101110001100;
        11'd1540: TDATA = 46'b0010010000110100010111001001101100001110111110;
        11'd1541: TDATA = 46'b0010010000011111100001101001101010101111110111;
        11'd1542: TDATA = 46'b0010010000001010101100101001101001010000110011;
        11'd1543: TDATA = 46'b0010001111110101111000001001100111110001110100;
        11'd1544: TDATA = 46'b0010001111100001000101001001100110010010111101;
        11'd1545: TDATA = 46'b0010001111001100010010101001100100110100001010;
        11'd1546: TDATA = 46'b0010001110110111100000001001100011010101011000;
        11'd1547: TDATA = 46'b0010001110100010101110101001100001110110101101;
        11'd1548: TDATA = 46'b0010001110001101111110001001100000011000001000;
        11'd1549: TDATA = 46'b0010001101111001001110001001011110111001100111;
        11'd1550: TDATA = 46'b0010001101100100011111101001011101011011001111;
        11'd1551: TDATA = 46'b0010001101001111110001001001011011111100111000;
        11'd1552: TDATA = 46'b0010001100111011000011001001011010011110100101;
        11'd1553: TDATA = 46'b0010001100100110010110001001011001000000011001;
        11'd1554: TDATA = 46'b0010001100010001101010001001010111100010010011;
        11'd1555: TDATA = 46'b0010001011111100111111001001010110000100010010;
        11'd1556: TDATA = 46'b0010001011101000010100101001010100100110010110;
        11'd1557: TDATA = 46'b0010001011010011101010001001010011001000011100;
        11'd1558: TDATA = 46'b0010001010111111000001101001010001101010101100;
        11'd1559: TDATA = 46'b0010001010101010011000101001010000001100111100;
        11'd1560: TDATA = 46'b0010001010010101110001001001001110101111010100;
        11'd1561: TDATA = 46'b0010001010000001001001101001001101010001101110;
        11'd1562: TDATA = 46'b0010001001101100100011101001001011110100010000;
        11'd1563: TDATA = 46'b0010001001010111111110001001001010010110110110;
        11'd1564: TDATA = 46'b0010001001000011011001001001001000111001100000;
        11'd1565: TDATA = 46'b0010001000101110110101001001000111011100010000;
        11'd1566: TDATA = 46'b0010001000011010010001101001000101111111000101;
        11'd1567: TDATA = 46'b0010001000000101101111101001000100100010000001;
        11'd1568: TDATA = 46'b0010000111110001001101001001000011000100111101;
        11'd1569: TDATA = 46'b0010000111011100101100001001000001101000000010;
        11'd1570: TDATA = 46'b0010000111001000001011101001000000001011001010;
        11'd1571: TDATA = 46'b0010000110110011101011101000111110101110010110;
        11'd1572: TDATA = 46'b0010000110011111001101001000111101010001101011;
        11'd1573: TDATA = 46'b0010000110001010101111001000111011110101000100;
        11'd1574: TDATA = 46'b0010000101110110010001001000111010011000011110;
        11'd1575: TDATA = 46'b0010000101100001110100101000111000111100000001;
        11'd1576: TDATA = 46'b0010000101001101011000101000110111011111100111;
        11'd1577: TDATA = 46'b0010000100111000111100101000110110000011010000;
        11'd1578: TDATA = 46'b0010000100100100100010001000110100100111000000;
        11'd1579: TDATA = 46'b0010000100010000001000001000110011001010110101;
        11'd1580: TDATA = 46'b0010000011111011101111001000110001101110101111;
        11'd1581: TDATA = 46'b0010000011100111010110101000110000010010101110;
        11'd1582: TDATA = 46'b0010000011010010111110101000101110110110110000;
        11'd1583: TDATA = 46'b0010000010111110100111101000101101011010111001;
        11'd1584: TDATA = 46'b0010000010101010010001001000101011111111000101;
        11'd1585: TDATA = 46'b0010000010010101111011101000101010100011011000;
        11'd1586: TDATA = 46'b0010000010000001100111001000101001000111110000;
        11'd1587: TDATA = 46'b0010000001101101010011001000100111101100001101;
        11'd1588: TDATA = 46'b0010000001011000111111001000100110010000101011;
        11'd1589: TDATA = 46'b0010000001000100101100001000100100110101001111;
        11'd1590: TDATA = 46'b0010000000110000011010101000100011011001111100;
        11'd1591: TDATA = 46'b0010000000011100001000101000100001111110101000;
        11'd1592: TDATA = 46'b0010000000000111111000001000100000100011011100;
        11'd1593: TDATA = 46'b0001111111110011101000001000011111001000010100;
        11'd1594: TDATA = 46'b0001111111011111011001001000011101101101010011;
        11'd1595: TDATA = 46'b0001111111001011001010101000011100010010010101;
        11'd1596: TDATA = 46'b0001111110110110111101001000011010110111011101;
        11'd1597: TDATA = 46'b0001111110100010101111101000011001011100100111;
        11'd1598: TDATA = 46'b0001111110001110100011001000011000000001110111;
        11'd1599: TDATA = 46'b0001111101111010010111101000010110100111001101;
        11'd1600: TDATA = 46'b0001111101100110001100101000010101001100100110;
        11'd1601: TDATA = 46'b0001111101010010000010001000010011110010000100;
        11'd1602: TDATA = 46'b0001111100111101111001001000010010010111101010;
        11'd1603: TDATA = 46'b0001111100101001110000001000010000111101010010;
        11'd1604: TDATA = 46'b0001111100010101101000001000001111100010111111;
        11'd1605: TDATA = 46'b0001111100000001100000101000001110001000110001;
        11'd1606: TDATA = 46'b0001111011101101011001101000001100101110100110;
        11'd1607: TDATA = 46'b0001111011011001010100001000001011010100100100;
        11'd1608: TDATA = 46'b0001111011000101001110101000001001111010100011;
        11'd1609: TDATA = 46'b0001111010110001001001101000001000100000100110;
        11'd1610: TDATA = 46'b0001111010011101000101101000000111000110101111;
        11'd1611: TDATA = 46'b0001111010001001000011001000000101101101000000;
        11'd1612: TDATA = 46'b0001111001110101000000101000000100010011010011;
        11'd1613: TDATA = 46'b0001111001100000111110101000000010111001101010;
        11'd1614: TDATA = 46'b0001111001001100111101001000000001100000000100;
        11'd1615: TDATA = 46'b0001111000111000111100101000000000000110100101;
        11'd1616: TDATA = 46'b0001111000100100111101000111111110101101001011;
        11'd1617: TDATA = 46'b0001111000010000111110000111111101010011110110;
        11'd1618: TDATA = 46'b0001110111111100111111100111111011111010100100;
        11'd1619: TDATA = 46'b0001110111101001000010100111111010100001011010;
        11'd1620: TDATA = 46'b0001110111010101000101000111111001001000010000;
        11'd1621: TDATA = 46'b0001110111000001001001000111110111101111001110;
        11'd1622: TDATA = 46'b0001110110101101001101100111110110010110010000;
        11'd1623: TDATA = 46'b0001110110011001010011000111110100111101011000;
        11'd1624: TDATA = 46'b0001110110000101011000100111110011100100100001;
        11'd1625: TDATA = 46'b0001110101110001011111000111110010001011110000;
        11'd1626: TDATA = 46'b0001110101011101100110100111110000110011000110;
        11'd1627: TDATA = 46'b0001110101001001101110100111101111011010011111;
        11'd1628: TDATA = 46'b0001110100110101110111000111101110000001111100;
        11'd1629: TDATA = 46'b0001110100100010000000100111101100101001011110;
        11'd1630: TDATA = 46'b0001110100001110001010100111101011010001000101;
        11'd1631: TDATA = 46'b0001110011111010010101000111101001111000110000;
        11'd1632: TDATA = 46'b0001110011100110100000100111101000100000100000;
        11'd1633: TDATA = 46'b0001110011010010101101000111100111001000010110;
        11'd1634: TDATA = 46'b0001110010111110111001100111100101110000001110;
        11'd1635: TDATA = 46'b0001110010101011000110100111100100011000001010;
        11'd1636: TDATA = 46'b0001110010010111010101000111100011000000001110;
        11'd1637: TDATA = 46'b0001110010000011100100000111100001101000010110;
        11'd1638: TDATA = 46'b0001110001101111110011100111100000010000100001;
        11'd1639: TDATA = 46'b0001110001011100000011100111011110111000110000;
        11'd1640: TDATA = 46'b0001110001001000010100100111011101100001000101;
        11'd1641: TDATA = 46'b0001110000110100100110100111011100001001100000;
        11'd1642: TDATA = 46'b0001110000100000111000100111011010110001111101;
        11'd1643: TDATA = 46'b0001110000001101001011000111011001011010011101;
        11'd1644: TDATA = 46'b0001101111111001011111000111011000000011000110;
        11'd1645: TDATA = 46'b0001101111100101110011000111010110101011110000;
        11'd1646: TDATA = 46'b0001101111010010001000100111010101010100100010;
        11'd1647: TDATA = 46'b0001101110111110011110000111010011111101010110;
        11'd1648: TDATA = 46'b0001101110101010110100100111010010100110001111;
        11'd1649: TDATA = 46'b0001101110010111001011100111010001001111001100;
        11'd1650: TDATA = 46'b0001101110000011100011000111001111111000001110;
        11'd1651: TDATA = 46'b0001101101101111111011100111001110100001010101;
        11'd1652: TDATA = 46'b0001101101011100010100100111001101001010011111;
        11'd1653: TDATA = 46'b0001101101001000101110100111001011110011110000;
        11'd1654: TDATA = 46'b0001101100110101001000100111001010011101000010;
        11'd1655: TDATA = 46'b0001101100100001100011100111001001000110011010;
        11'd1656: TDATA = 46'b0001101100001101111111100111000111101111111000;
        11'd1657: TDATA = 46'b0001101011111010011100000111000110011001011010;
        11'd1658: TDATA = 46'b0001101011100110111001000111000101000010111111;
        11'd1659: TDATA = 46'b0001101011010011010111100111000011101100101101;
        11'd1660: TDATA = 46'b0001101010111111110101100111000010010110011010;
        11'd1661: TDATA = 46'b0001101010101100010100100111000001000000001100;
        11'd1662: TDATA = 46'b0001101010011000110100100110111111101010000101;
        11'd1663: TDATA = 46'b0001101010000101010101000110111110010100000001;
        11'd1664: TDATA = 46'b0001101001110001110110100110111100111110000011;
        11'd1665: TDATA = 46'b0001101001011110011000000110111011101000000111;
        11'd1666: TDATA = 46'b0001101001001010111011000110111010010010010011;
        11'd1667: TDATA = 46'b0001101000110111011101100110111000111100011110;
        11'd1668: TDATA = 46'b0001101000100100000001000110110111100110101111;
        11'd1669: TDATA = 46'b0001101000010000100110100110110110010001001010;
        11'd1670: TDATA = 46'b0001100111111101001011100110110100111011100101;
        11'd1671: TDATA = 46'b0001100111101001110001000110110011100110000011;
        11'd1672: TDATA = 46'b0001100111010110010111100110110010010000100111;
        11'd1673: TDATA = 46'b0001100111000010111111000110110000111011010001;
        11'd1674: TDATA = 46'b0001100110101111100111000110101111100101111110;
        11'd1675: TDATA = 46'b0001100110011100001111100110101110010000110000;
        11'd1676: TDATA = 46'b0001100110001000111000100110101100111011100101;
        11'd1677: TDATA = 46'b0001100101110101100010100110101011100110011111;
        11'd1678: TDATA = 46'b0001100101100010001101000110101010010001011110;
        11'd1679: TDATA = 46'b0001100101001110111000000110101000111100100000;
        11'd1680: TDATA = 46'b0001100100111011100100000110100111100111101000;
        11'd1681: TDATA = 46'b0001100100101000010001000110100110010010110110;
        11'd1682: TDATA = 46'b0001100100010100111101100110100100111110000011;
        11'd1683: TDATA = 46'b0001100100000001101011100110100011101001011000;
        11'd1684: TDATA = 46'b0001100011101110011010000110100010010100110001;
        11'd1685: TDATA = 46'b0001100011011011001001000110100001000000001101;
        11'd1686: TDATA = 46'b0001100011000111111001000110011111101011101111;
        11'd1687: TDATA = 46'b0001100010110100101001100110011110010111010101;
        11'd1688: TDATA = 46'b0001100010100001011010100110011101000010111111;
        11'd1689: TDATA = 46'b0001100010001110001100100110011011101110101110;
        11'd1690: TDATA = 46'b0001100001111010111111000110011010011010100001;
        11'd1691: TDATA = 46'b0001100001100111110010000110011001000110011000;
        11'd1692: TDATA = 46'b0001100001010100100110000110010111110010010100;
        11'd1693: TDATA = 46'b0001100001000001011010100110010110011110010100;
        11'd1694: TDATA = 46'b0001100000101110001111100110010101001010011000;
        11'd1695: TDATA = 46'b0001100000011011000101000110010011110110011111;
        11'd1696: TDATA = 46'b0001100000000111111011100110010010100010101100;
        11'd1697: TDATA = 46'b0001011111110100110010100110010001001110111101;
        11'd1698: TDATA = 46'b0001011111100001101010100110001111111011010100;
        11'd1699: TDATA = 46'b0001011111001110100011000110001110100111101110;
        11'd1700: TDATA = 46'b0001011110111011011100000110001101010100001100;
        11'd1701: TDATA = 46'b0001011110101000010101000110001100000000101011;
        11'd1702: TDATA = 46'b0001011110010101001111100110001010101101010010;
        11'd1703: TDATA = 46'b0001011110000010001011000110001001011001111111;
        11'd1704: TDATA = 46'b0001011101101111000111000110001000000110110000;
        11'd1705: TDATA = 46'b0001011101011100000011000110000110110011100010;
        11'd1706: TDATA = 46'b0001011101001000111111100110000101100000010111;
        11'd1707: TDATA = 46'b0001011100110101111101000110000100001101010011;
        11'd1708: TDATA = 46'b0001011100100010111100000110000010111010010110;
        11'd1709: TDATA = 46'b0001011100001111111010000110000001100111010110;
        11'd1710: TDATA = 46'b0001011011111100111010000110000000010100100001;
        11'd1711: TDATA = 46'b0001011011101001111010000101111111000001101101;
        11'd1712: TDATA = 46'b0001011011010110111011000101111101101110111110;
        11'd1713: TDATA = 46'b0001011011000011111100000101111100011100010010;
        11'd1714: TDATA = 46'b0001011010110000111110100101111011001001101101;
        11'd1715: TDATA = 46'b0001011010011110000001000101111001110111001001;
        11'd1716: TDATA = 46'b0001011010001011000100100101111000100100101011;
        11'd1717: TDATA = 46'b0001011001111000001000100101110111010010010001;
        11'd1718: TDATA = 46'b0001011001100101001101000101110101111111111010;
        11'd1719: TDATA = 46'b0001011001010010010010100101110100101101101010;
        11'd1720: TDATA = 46'b0001011000111111011000000101110011011011011010;
        11'd1721: TDATA = 46'b0001011000101100011111000101110010001001010011;
        11'd1722: TDATA = 46'b0001011000011001100110100101110000110111001111;
        11'd1723: TDATA = 46'b0001011000000110101101100101101111100101001010;
        11'd1724: TDATA = 46'b0001010111110011110110100101101110010011001111;
        11'd1725: TDATA = 46'b0001010111100000111111100101101101000001010110;
        11'd1726: TDATA = 46'b0001010111001110001010000101101011101111100100;
        11'd1727: TDATA = 46'b0001010110111011010100000101101010011101110010;
        11'd1728: TDATA = 46'b0001010110101000011111000101101001001100000110;
        11'd1729: TDATA = 46'b0001010110010101101011000101100111111010011111;
        11'd1730: TDATA = 46'b0001010110000010110111000101100110101000111001;
        11'd1731: TDATA = 46'b0001010101110000000100000101100101010111011010;
        11'd1732: TDATA = 46'b0001010101011101010001100101100100000101111110;
        11'd1733: TDATA = 46'b0001010101001010100000100101100010110100101010;
        11'd1734: TDATA = 46'b0001010100110111101111000101100001100011010100;
        11'd1735: TDATA = 46'b0001010100100100111110100101100000010010000101;
        11'd1736: TDATA = 46'b0001010100010010001111000101011111000000111100;
        11'd1737: TDATA = 46'b0001010011111111011111100101011101101111110011;
        11'd1738: TDATA = 46'b0001010011101100110001100101011100011110110011;
        11'd1739: TDATA = 46'b0001010011011010000011000101011011001101110010;
        11'd1740: TDATA = 46'b0001010011000111010101100101011001111100110110;
        11'd1741: TDATA = 46'b0001010010110100101001000101011000101100000001;
        11'd1742: TDATA = 46'b0001010010100001111101000101010111011011001110;
        11'd1743: TDATA = 46'b0001010010001111010001100101010110001010100000;
        11'd1744: TDATA = 46'b0001010001111100100111000101010100111001110111;
        11'd1745: TDATA = 46'b0001010001101001111101000101010011101001010001;
        11'd1746: TDATA = 46'b0001010001010111010011100101010010011000101111;
        11'd1747: TDATA = 46'b0001010001000100101010100101010001001000010000;
        11'd1748: TDATA = 46'b0001010000110010000010100101001111110111111000;
        11'd1749: TDATA = 46'b0001010000011111011010100101001110100111100000;
        11'd1750: TDATA = 46'b0001010000001100110011100101001101010111001110;
        11'd1751: TDATA = 46'b0001001111111010001101000101001100000111000000;
        11'd1752: TDATA = 46'b0001001111100111100111100101001010110110111000;
        11'd1753: TDATA = 46'b0001001111010101000010100101001001100110110010;
        11'd1754: TDATA = 46'b0001001111000010011101100101001000010110101111;
        11'd1755: TDATA = 46'b0001001110101111111001100101000111000110110001;
        11'd1756: TDATA = 46'b0001001110011101010111000101000101110110111010;
        11'd1757: TDATA = 46'b0001001110001010110100100101000100100111000101;
        11'd1758: TDATA = 46'b0001001101111000010010100101000011010111010100;
        11'd1759: TDATA = 46'b0001001101100101110000100101000010000111100100;
        11'd1760: TDATA = 46'b0001001101010011010000000101000000110111111011;
        11'd1761: TDATA = 46'b0001001101000000110000000100111111101000010110;
        11'd1762: TDATA = 46'b0001001100101110010000000100111110011000110011;
        11'd1763: TDATA = 46'b0001001100011011110001100100111101001001010111;
        11'd1764: TDATA = 46'b0001001100001001010011100100111011111001111111;
        11'd1765: TDATA = 46'b0001001011110110110101100100111010101010101000;
        11'd1766: TDATA = 46'b0001001011100100011000100100111001011011010111;
        11'd1767: TDATA = 46'b0001001011010001111100100100111000001100001011;
        11'd1768: TDATA = 46'b0001001010111111100000100100110110111101000001;
        11'd1769: TDATA = 46'b0001001010101101000101000100110101101101111010;
        11'd1770: TDATA = 46'b0001001010011010101011000100110100011110111011;
        11'd1771: TDATA = 46'b0001001010001000010000100100110011001111111011;
        11'd1772: TDATA = 46'b0001001001110101110111000100110010000001000001;
        11'd1773: TDATA = 46'b0001001001100011011110100100110000110010001100;
        11'd1774: TDATA = 46'b0001001001010001000110100100101111100011011011;
        11'd1775: TDATA = 46'b0001001000111110101111000100101110010100101101;
        11'd1776: TDATA = 46'b0001001000101100011000100100101101000110000101;
        11'd1777: TDATA = 46'b0001001000011010000010000100101011110111011110;
        11'd1778: TDATA = 46'b0001001000000111101100100100101010101000111101;
        11'd1779: TDATA = 46'b0001000111110101010111100100101001011010011111;
        11'd1780: TDATA = 46'b0001000111100011000011000100101000001100000100;
        11'd1781: TDATA = 46'b0001000111010000101111000100100110111101101110;
        11'd1782: TDATA = 46'b0001000110111110011100000100100101101111011100;
        11'd1783: TDATA = 46'b0001000110101100001001100100100100100001001110;
        11'd1784: TDATA = 46'b0001000110011001110111100100100011010011000100;
        11'd1785: TDATA = 46'b0001000110000111100110100100100010000100111111;
        11'd1786: TDATA = 46'b0001000101110101010101100100100000110110111100;
        11'd1787: TDATA = 46'b0001000101100011000101100100011111101000111110;
        11'd1788: TDATA = 46'b0001000101010000110101100100011110011011000001;
        11'd1789: TDATA = 46'b0001000100111110100111000100011101001101001100;
        11'd1790: TDATA = 46'b0001000100101100011000100100011011111111011000;
        11'd1791: TDATA = 46'b0001000100011010001010100100011010110001101000;
        11'd1792: TDATA = 46'b0001000100000111111101100100011001100011111101;
        11'd1793: TDATA = 46'b0001000011110101110001000100011000010110010110;
        11'd1794: TDATA = 46'b0001000011100011100101000100010111001000110010;
        11'd1795: TDATA = 46'b0001000011010001011010100100010101111011010110;
        11'd1796: TDATA = 46'b0001000010111111001111100100010100101101111001;
        11'd1797: TDATA = 46'b0001000010101101000101100100010011100000100010;
        11'd1798: TDATA = 46'b0001000010011010111100100100010010010011010000;
        11'd1799: TDATA = 46'b0001000010001000110011100100010001000101111111;
        11'd1800: TDATA = 46'b0001000001110110101011000100001111111000110010;
        11'd1801: TDATA = 46'b0001000001100100100011000100001110101011101000;
        11'd1802: TDATA = 46'b0001000001010010011100100100001101011110100110;
        11'd1803: TDATA = 46'b0001000001000000010101100100001100010001100011;
        11'd1804: TDATA = 46'b0001000000101110010000000100001011000100101000;
        11'd1805: TDATA = 46'b0001000000011100001011000100001001110111110000;
        11'd1806: TDATA = 46'b0001000000001010000110100100001000101010111100;
        11'd1807: TDATA = 46'b0000111111111000000001100100000111011110000110;
        11'd1808: TDATA = 46'b0000111111100101111111000100000110010001011101;
        11'd1809: TDATA = 46'b0000111111010011111100000100000101000100110011;
        11'd1810: TDATA = 46'b0000111111000001111001100100000011111000001100;
        11'd1811: TDATA = 46'b0000111110101111111000000100000010101011101011;
        11'd1812: TDATA = 46'b0000111110011101110111000100000001011111001101;
        11'd1813: TDATA = 46'b0000111110001011110110100100000000010010110010;
        11'd1814: TDATA = 46'b0000111101111001110110100011111111000110011011;
        11'd1815: TDATA = 46'b0000111101100111110111100011111101111010001001;
        11'd1816: TDATA = 46'b0000111101010101111000100011111100101101111001;
        11'd1817: TDATA = 46'b0000111101000011111011000011111011100001110000;
        11'd1818: TDATA = 46'b0000111100110001111101000011111010010101100110;
        11'd1819: TDATA = 46'b0000111100100000000000100011111001001001100100;
        11'd1820: TDATA = 46'b0000111100001110000100100011110111111101100101;
        11'd1821: TDATA = 46'b0000111011111100001000100011110110110001101000;
        11'd1822: TDATA = 46'b0000111011101010001101000011110101100101101110;
        11'd1823: TDATA = 46'b0000111011011000010011000011110100011001111100;
        11'd1824: TDATA = 46'b0000111011000110011001000011110011001110001010;
        11'd1825: TDATA = 46'b0000111010110100011111100011110010000010011101;
        11'd1826: TDATA = 46'b0000111010100010100111000011110000110110110100;
        11'd1827: TDATA = 46'b0000111010010000101110100011101111101011001101;
        11'd1828: TDATA = 46'b0000111001111110110111000011101110011111101011;
        11'd1829: TDATA = 46'b0000111001101101000000000011101101010100001101;
        11'd1830: TDATA = 46'b0000111001011011001010000011101100001000110100;
        11'd1831: TDATA = 46'b0000111001001001010100000011101010111101011101;
        11'd1832: TDATA = 46'b0000111000110111011111000011101001110010001011;
        11'd1833: TDATA = 46'b0000111000100101101010000011101000100110111010;
        11'd1834: TDATA = 46'b0000111000010011110110100011100111011011110001;
        11'd1835: TDATA = 46'b0000111000000010000011000011100110010000101001;
        11'd1836: TDATA = 46'b0000110111110000010000000011100101000101100100;
        11'd1837: TDATA = 46'b0000110111011110011101100011100011111010100011;
        11'd1838: TDATA = 46'b0000110111001100101100000011100010101111100111;
        11'd1839: TDATA = 46'b0000110110111010111011000011100001100100101110;
        11'd1840: TDATA = 46'b0000110110101001001010100011100000011001111001;
        11'd1841: TDATA = 46'b0000110110010111011010100011011111001111000111;
        11'd1842: TDATA = 46'b0000110110000101101011100011011110000100011011;
        11'd1843: TDATA = 46'b0000110101110011111100100011011100111001110000;
        11'd1844: TDATA = 46'b0000110101100010001110100011011011101111001010;
        11'd1845: TDATA = 46'b0000110101010000100001000011011010100100100111;
        11'd1846: TDATA = 46'b0000110100111110110100000011011001011010001000;
        11'd1847: TDATA = 46'b0000110100101101000111100011011000001111101100;
        11'd1848: TDATA = 46'b0000110100011011011011100011010111000101010100;
        11'd1849: TDATA = 46'b0000110100001001110000100011010101111011000001;
        11'd1850: TDATA = 46'b0000110011111000000101100011010100110000101111;
        11'd1851: TDATA = 46'b0000110011100110011011100011010011100110100011;
        11'd1852: TDATA = 46'b0000110011010100110010000011010010011100011010;
        11'd1853: TDATA = 46'b0000110011000011001001100011010001010010010110;
        11'd1854: TDATA = 46'b0000110010110001100000100011010000001000010010;
        11'd1855: TDATA = 46'b0000110010011111111001000011001110111110010101;
        11'd1856: TDATA = 46'b0000110010001110010001100011001101110100011001;
        11'd1857: TDATA = 46'b0000110001111100101011000011001100101010100010;
        11'd1858: TDATA = 46'b0000110001101011000101000011001011100000101111;
        11'd1859: TDATA = 46'b0000110001011001011111100011001010010111000000;
        11'd1860: TDATA = 46'b0000110001000111111011000011001001001101010101;
        11'd1861: TDATA = 46'b0000110000110110010111000011001000000011101110;
        11'd1862: TDATA = 46'b0000110000100100110011000011000110111010001000;
        11'd1863: TDATA = 46'b0000110000010011001111100011000101110000100110;
        11'd1864: TDATA = 46'b0000110000000001101101000011000100100111001000;
        11'd1865: TDATA = 46'b0000101111110000001010100011000011011101101100;
        11'd1866: TDATA = 46'b0000101111011110101001100011000010010100011000;
        11'd1867: TDATA = 46'b0000101111001101001000100011000001001011000101;
        11'd1868: TDATA = 46'b0000101110111011101000000011000000000001110101;
        11'd1869: TDATA = 46'b0000101110101010001000100010111110111000101010;
        11'd1870: TDATA = 46'b0000101110011000101001100010111101101111100011;
        11'd1871: TDATA = 46'b0000101110000111001011000010111100100110011111;
        11'd1872: TDATA = 46'b0000101101110101101100100010111011011101011100;
        11'd1873: TDATA = 46'b0000101101100100001111100010111010010100100000;
        11'd1874: TDATA = 46'b0000101101010010110010100010111001001011100110;
        11'd1875: TDATA = 46'b0000101101000001010110100010111000000010110001;
        11'd1876: TDATA = 46'b0000101100101111111010100010110110111001111110;
        11'd1877: TDATA = 46'b0000101100011110011111000010110101110001001101;
        11'd1878: TDATA = 46'b0000101100001101000100100010110100101000100010;
        11'd1879: TDATA = 46'b0000101011111011101011000010110011011111111100;
        11'd1880: TDATA = 46'b0000101011101010010001000010110010010111010110;
        11'd1881: TDATA = 46'b0000101011011000111000000010110001001110110101;
        11'd1882: TDATA = 46'b0000101011000111100000000010110000000110011001;
        11'd1883: TDATA = 46'b0000101010110110001000100010101110111110000000;
        11'd1884: TDATA = 46'b0000101010100100110000100010101101110101100111;
        11'd1885: TDATA = 46'b0000101010010011011010100010101100101101010111;
        11'd1886: TDATA = 46'b0000101010000010000100000010101011100101000110;
        11'd1887: TDATA = 46'b0000101001110000101111000010101010011100111100;
        11'd1888: TDATA = 46'b0000101001011111011001100010101001010100110010;
        11'd1889: TDATA = 46'b0000101001001110000101100010101000001100101111;
        11'd1890: TDATA = 46'b0000101000111100110001100010100111000100101101;
        11'd1891: TDATA = 46'b0000101000101011011110100010100101111100110000;
        11'd1892: TDATA = 46'b0000101000011010001011100010100100110100110101;
        11'd1893: TDATA = 46'b0000101000001000111001100010100011101100111111;
        11'd1894: TDATA = 46'b0000100111110111101000000010100010100101001100;
        11'd1895: TDATA = 46'b0000100111100110010110100010100001011101011011;
        11'd1896: TDATA = 46'b0000100111010101000110100010100000010101110001;
        11'd1897: TDATA = 46'b0000100111000011110110100010011111001110001000;
        11'd1898: TDATA = 46'b0000100110110010100111100010011110000110100100;
        11'd1899: TDATA = 46'b0000100110100001011000100010011100111111000001;
        11'd1900: TDATA = 46'b0000100110010000001010100010011011110111100100;
        11'd1901: TDATA = 46'b0000100101111110111101000010011010110000001010;
        11'd1902: TDATA = 46'b0000100101101101101111100010011001101000110001;
        11'd1903: TDATA = 46'b0000100101011100100011000010011000100001011110;
        11'd1904: TDATA = 46'b0000100101001011010111000010010111011010001101;
        11'd1905: TDATA = 46'b0000100100111010001011100010010110010011000000;
        11'd1906: TDATA = 46'b0000100100101001000000100010010101001011110110;
        11'd1907: TDATA = 46'b0000100100010111110110000010010100000100110000;
        11'd1908: TDATA = 46'b0000100100000110101100100010010010111101101110;
        11'd1909: TDATA = 46'b0000100011110101100011100010010001110110110000;
        11'd1910: TDATA = 46'b0000100011100100011011000010010000101111110101;
        11'd1911: TDATA = 46'b0000100011010011010010100010001111101000111100;
        11'd1912: TDATA = 46'b0000100011000010001011000010001110100010000111;
        11'd1913: TDATA = 46'b0000100010110001000100000010001101011011010110;
        11'd1914: TDATA = 46'b0000100010011111111101100010001100010100101000;
        11'd1915: TDATA = 46'b0000100010001110111000000010001011001101111111;
        11'd1916: TDATA = 46'b0000100001111101110010100010001010000111010111;
        11'd1917: TDATA = 46'b0000100001101100101101100010001001000000110011;
        11'd1918: TDATA = 46'b0000100001011011101001100010000111111010010100;
        11'd1919: TDATA = 46'b0000100001001010100101100010000110110011110110;
        11'd1920: TDATA = 46'b0000100000111001100010100010000101101101011101;
        11'd1921: TDATA = 46'b0000100000101000100000000010000100100111000111;
        11'd1922: TDATA = 46'b0000100000010111011110000010000011100000110101;
        11'd1923: TDATA = 46'b0000100000000110011100100010000010011010100110;
        11'd1924: TDATA = 46'b0000011111110101011100000010000001010100011100;
        11'd1925: TDATA = 46'b0000011111100100011011100010000000001110010011;
        11'd1926: TDATA = 46'b0000011111010011011011100001111111001000001101;
        11'd1927: TDATA = 46'b0000011111000010011100000001111110000010001011;
        11'd1928: TDATA = 46'b0000011110110001011101100001111100111100001110;
        11'd1929: TDATA = 46'b0000011110100000011111100001111011110110010100;
        11'd1930: TDATA = 46'b0000011110001111100001100001111010110000011011;
        11'd1931: TDATA = 46'b0000011101111110100100100001111001101010100111;
        11'd1932: TDATA = 46'b0000011101101101101000100001111000100100111001;
        11'd1933: TDATA = 46'b0000011101011100101100100001110111011111001100;
        11'd1934: TDATA = 46'b0000011101001011110000100001110110011001100000;
        11'd1935: TDATA = 46'b0000011100111010110101100001110101010011111001;
        11'd1936: TDATA = 46'b0000011100101001111011000001110100001110010101;
        11'd1937: TDATA = 46'b0000011100011001000001000001110011001000110100;
        11'd1938: TDATA = 46'b0000011100001000001000000001110010000011011001;
        11'd1939: TDATA = 46'b0000011011110111001111000001110000111101111111;
        11'd1940: TDATA = 46'b0000011011100110010111000001101111111000101010;
        11'd1941: TDATA = 46'b0000011011010101011111000001101110110011010110;
        11'd1942: TDATA = 46'b0000011011000100101000000001101101101110000111;
        11'd1943: TDATA = 46'b0000011010110011110001100001101100101000111100;
        11'd1944: TDATA = 46'b0000011010100010111011100001101011100011110011;
        11'd1945: TDATA = 46'b0000011010010010000110000001101010011110101110;
        11'd1946: TDATA = 46'b0000011010000001010001000001101001011001101100;
        11'd1947: TDATA = 46'b0000011001110000011100100001101000010100101101;
        11'd1948: TDATA = 46'b0000011001011111101001000001100111001111110100;
        11'd1949: TDATA = 46'b0000011001001110110101100001100110001010111011;
        11'd1950: TDATA = 46'b0000011000111110000010100001100101000110000110;
        11'd1951: TDATA = 46'b0000011000101101010000100001100100000001010110;
        11'd1952: TDATA = 46'b0000011000011100011110100001100010111100100110;
        11'd1953: TDATA = 46'b0000011000001011101101000001100001110111111010;
        11'd1954: TDATA = 46'b0000010111111010111100100001100000110011010100;
        11'd1955: TDATA = 46'b0000010111101010001100100001011111101110110000;
        11'd1956: TDATA = 46'b0000010111011001011101000001011110101010010000;
        11'd1957: TDATA = 46'b0000010111001000101101100001011101100101110000;
        11'd1958: TDATA = 46'b0000010110110111111111100001011100100001011000;
        11'd1959: TDATA = 46'b0000010110100111010001100001011011011101000001;
        11'd1960: TDATA = 46'b0000010110010110100100000001011010011000101101;
        11'd1961: TDATA = 46'b0000010110000101110111000001011001010100011100;
        11'd1962: TDATA = 46'b0000010101110101001010100001011000010000001111;
        11'd1963: TDATA = 46'b0000010101100100011110100001010111001100000100;
        11'd1964: TDATA = 46'b0000010101010011110011100001010110000111111111;
        11'd1965: TDATA = 46'b0000010101000011001000100001010101000011111010;
        11'd1966: TDATA = 46'b0000010100110010011110000001010011111111111001;
        11'd1967: TDATA = 46'b0000010100100001110100100001010010111011111101;
        11'd1968: TDATA = 46'b0000010100010001001011100001010001111000000100;
        11'd1969: TDATA = 46'b0000010100000000100010100001010000110100001101;
        11'd1970: TDATA = 46'b0000010011101111111010100001001111110000011010;
        11'd1971: TDATA = 46'b0000010011011111010011000001001110101100101011;
        11'd1972: TDATA = 46'b0000010011001110101100000001001101101000111110;
        11'd1973: TDATA = 46'b0000010010111110000101000001001100100101010011;
        11'd1974: TDATA = 46'b0000010010101101011111000001001011100001101101;
        11'd1975: TDATA = 46'b0000010010011100111001100001001010011110001010;
        11'd1976: TDATA = 46'b0000010010001100010101000001001001011010101100;
        11'd1977: TDATA = 46'b0000010001111011110000100001001000010111001111;
        11'd1978: TDATA = 46'b0000010001101011001100100001000111010011110101;
        11'd1979: TDATA = 46'b0000010001011010101001000001000110010000011111;
        11'd1980: TDATA = 46'b0000010001001010000110100001000101001101001101;
        11'd1981: TDATA = 46'b0000010000111001100100000001000100001001111101;
        11'd1982: TDATA = 46'b0000010000101001000010000001000011000110101111;
        11'd1983: TDATA = 46'b0000010000011000100000100001000010000011100101;
        11'd1984: TDATA = 46'b0000010000001000000000000001000001000000100000;
        11'd1985: TDATA = 46'b0000001111110111011111100000111111111101011100;
        11'd1986: TDATA = 46'b0000001111100111000000000000111110111010011101;
        11'd1987: TDATA = 46'b0000001111010110100000100000111101110111011111;
        11'd1988: TDATA = 46'b0000001111000110000010000000111100110100100111;
        11'd1989: TDATA = 46'b0000001110110101100100000000111011110001110001;
        11'd1990: TDATA = 46'b0000001110100101000110100000111010101110111111;
        11'd1991: TDATA = 46'b0000001110010100101001000000111001101100001101;
        11'd1992: TDATA = 46'b0000001110000100001100100000111000101001100001;
        11'd1993: TDATA = 46'b0000001101110011110000100000110111100110110111;
        11'd1994: TDATA = 46'b0000001101100011010101000000110110100100010001;
        11'd1995: TDATA = 46'b0000001101010010111010000000110101100001101110;
        11'd1996: TDATA = 46'b0000001101000010011111100000110100011111001110;
        11'd1997: TDATA = 46'b0000001100110010000101100000110011011100110001;
        11'd1998: TDATA = 46'b0000001100100001101100000000110010011010010111;
        11'd1999: TDATA = 46'b0000001100010001010011000000110001011000000000;
        11'd2000: TDATA = 46'b0000001100000000111010100000110000010101101101;
        11'd2001: TDATA = 46'b0000001011110000100010100000101111010011011100;
        11'd2002: TDATA = 46'b0000001011100000001011100000101110010001010001;
        11'd2003: TDATA = 46'b0000001011001111110100100000101101001111000110;
        11'd2004: TDATA = 46'b0000001010111111011110000000101100001100111111;
        11'd2005: TDATA = 46'b0000001010101111001000100000101011001010111100;
        11'd2006: TDATA = 46'b0000001010011110110011000000101010001000111011;
        11'd2007: TDATA = 46'b0000001010001110011110000000101001000110111101;
        11'd2008: TDATA = 46'b0000001001111110001010000000101000000101000011;
        11'd2009: TDATA = 46'b0000001001101101110110100000100111000011001101;
        11'd2010: TDATA = 46'b0000001001011101100011000000100110000001011000;
        11'd2011: TDATA = 46'b0000001001001101010000000000100100111111100110;
        11'd2012: TDATA = 46'b0000001000111100111101100000100011111101110111;
        11'd2013: TDATA = 46'b0000001000101100101100100000100010111100001111;
        11'd2014: TDATA = 46'b0000001000011100011010100000100001111010100100;
        11'd2015: TDATA = 46'b0000001000001100001010000000100000111001000001;
        11'd2016: TDATA = 46'b0000000111111011111010000000011111110111100000;
        11'd2017: TDATA = 46'b0000000111101011101010000000011110110110000000;
        11'd2018: TDATA = 46'b0000000111011011011011100000011101110100100111;
        11'd2019: TDATA = 46'b0000000111001011001100100000011100110011001110;
        11'd2020: TDATA = 46'b0000000110111010111110100000011011110001111001;
        11'd2021: TDATA = 46'b0000000110101010110001000000011010110000101000;
        11'd2022: TDATA = 46'b0000000110011010100011100000011001101111010111;
        11'd2023: TDATA = 46'b0000000110001010010111000000011000101110001100;
        11'd2024: TDATA = 46'b0000000101111010001011000000010111101101000011;
        11'd2025: TDATA = 46'b0000000101101001111111100000010110101011111110;
        11'd2026: TDATA = 46'b0000000101011001110100100000010101101010111100;
        11'd2027: TDATA = 46'b0000000101001001101001100000010100101001111010;
        11'd2028: TDATA = 46'b0000000100111001011111100000010011101000111110;
        11'd2029: TDATA = 46'b0000000100101001010110000000010010101000000101;
        11'd2030: TDATA = 46'b0000000100011001001101000000010001100111001110;
        11'd2031: TDATA = 46'b0000000100001001000100100000010000100110011011;
        11'd2032: TDATA = 46'b0000000011111000111100100000001111100101101011;
        11'd2033: TDATA = 46'b0000000011101000110101000000001110100100111110;
        11'd2034: TDATA = 46'b0000000011011000101101100000001101100100010010;
        11'd2035: TDATA = 46'b0000000011001000100111000000001100100011101011;
        11'd2036: TDATA = 46'b0000000010111000100001000000001011100011000110;
        11'd2037: TDATA = 46'b0000000010101000011011100000001010100010100101;
        11'd2038: TDATA = 46'b0000000010011000010111000000001001100010001001;
        11'd2039: TDATA = 46'b0000000010001000010001100000001000100001101010;
        11'd2040: TDATA = 46'b0000000001111000001101100000000111100001010010;
        11'd2041: TDATA = 46'b0000000001101000001011000000000110100001000001;
        11'd2042: TDATA = 46'b0000000001011000000111100000000101100000101101;
        11'd2043: TDATA = 46'b0000000001001000000101000000000100100000011110;
        11'd2044: TDATA = 46'b0000000000111000000011100000000011100000010100;
        11'd2045: TDATA = 46'b0000000000101000000001100000000010100000001001;
        11'd2046: TDATA = 46'b0000000000011000000000100000000001100000000011;
        11'd2047: TDATA = 46'b0000000000001000000000000000000000100000000000;
	endcase
    end
    endfunction

    assign tdata = TDATA(mal);
    
    wire [22:0] mx0,mx02;
    assign mx0 = tdata[45:23];
    assign mx02 = tdata[22:0];

    wire [47:0] max02a;
    assign max02a = {1'b1,ma} * {1'b1,mx02};

    wire [22:0] max02;
    assign max02 = (max02a[47:47]) ? max02a[46:24]: max02a[45:23];

    wire [24:0] mix2a;
    assign mix2a = {1'b1,mx0,1'b0} - {2'b01,max02};

    wire [22:0] mix2;
    assign mix2 = mix2a[22:0];

    wire six2;
    assign six2 = sa;

    wire [7:0] eb;
    assign eb = 8'd253;

    wire sx,sy;
    wire [7:0] ex,ey;
    wire [22:0] mx,my;
    assign sx = x1[31:31];
    assign ex = x1[30:23];
    assign mx = x1[22:0];

    assign sy = sx ^ six2;

    wire [47:0] mya;
    assign mya = {1'b1,mx} * {1'b1,mix2};

    wire a;
    assign a = mya[47:47];
    assign my = (a) ? mya[46:24]: mya[45:23];

    wire [7:0] e2ab;
    assign e2ab = (ex == 8'b0) ? 0: eb;

    wire [8:0] eya;
    assign eya = ex + e2ab + a;

    wire [8:0] eyb;
    assign eyb = 9'd127 + ea;

    assign ey = (eya > eyb) ? eya - eyb: 0;

    assign y = {sy,ey,my};

endmodule
