
module fsqrt(
    input wire [31:0] x,
    output wire [31:0] y);

    wire odd_flag;
    wire [7:0] ex;
    wire [22:0] mx;
    wire [11:0] index;
    assign odd_flag = x[23:23];
    assign ex = x[30:23];
    assign mx = x[22:0];
    assign index = x[23:12];

    function [49:0] TDATA (
	input [11:0] INDEX
    );
    begin
	casex(INDEX)
        12'd0: TDATA = 50'b10000111101111110111100011011010011110011111110110;
        12'd1: TDATA = 50'b10000111101101101111111001011010011010010000101011;
        12'd2: TDATA = 50'b10000111101011101000010101011010010110000001110100;
        12'd3: TDATA = 50'b10000111101001100000110111011010010001110011010001;
        12'd4: TDATA = 50'b10000111100111011001100001011010001101100101001001;
        12'd5: TDATA = 50'b10000111100101010010001101011010001001010111001001;
        12'd6: TDATA = 50'b10000111100011001011000011011010000101001001101001;
        12'd7: TDATA = 50'b10000111100001000100000011011010000000111100100100;
        12'd8: TDATA = 50'b10000111011110111101000001011001111100101111100001;
        12'd9: TDATA = 50'b10000111011100110110001001011001111000100010111111;
        12'd10: TDATA = 50'b10000111011010101111011001011001110100010110110001;
        12'd11: TDATA = 50'b10000111011000101000101011011001110000001010110001;
        12'd12: TDATA = 50'b10000111010110100010000011011001101011111111000101;
        12'd13: TDATA = 50'b10000111010100011011100111011001100111110011111010;
        12'd14: TDATA = 50'b10000111010010010101010001011001100011101001000011;
        12'd15: TDATA = 50'b10000111010000001110111011011001011111011110010100;
        12'd16: TDATA = 50'b10000111001110001000110001011001011011010100000101;
        12'd17: TDATA = 50'b10000111001100000010101001011001010111001010000100;
        12'd18: TDATA = 50'b10000111001001111100101011011001010011000000011101;
        12'd19: TDATA = 50'b10000111000111110110110011011001001110110111001011;
        12'd20: TDATA = 50'b10000111000101110000111111011001001010101110000111;
        12'd21: TDATA = 50'b10000111000011101011010011011001000110100101011100;
        12'd22: TDATA = 50'b10000111000001100101101101011001000010011101000110;
        12'd23: TDATA = 50'b10000110111111100000001101011000111110010101000100;
        12'd24: TDATA = 50'b10000110111101011010101111011000111010001101010000;
        12'd25: TDATA = 50'b10000110111011010101011001011000110110000101110000;
        12'd26: TDATA = 50'b10000110111001010000001011011000110001111110101001;
        12'd27: TDATA = 50'b10000110110111001011000011011000101101110111110111;
        12'd28: TDATA = 50'b10000110110101000110000111011000101001110001100101;
        12'd29: TDATA = 50'b10000110110011000001000111011000100101101011010100;
        12'd30: TDATA = 50'b10000110110000111100010101011000100001100101100100;
        12'd31: TDATA = 50'b10000110101110110111100001011000011101011111111011;
        12'd32: TDATA = 50'b10000110101100110010111011011000011001011010110010;
        12'd33: TDATA = 50'b10000110101010101110010111011000010101010101110111;
        12'd34: TDATA = 50'b10000110101000101001111001011000010001010001010000;
        12'd35: TDATA = 50'b10000110100110100101100011011000001101001101000011;
        12'd36: TDATA = 50'b10000110100100100001010001011000001001001001000011;
        12'd37: TDATA = 50'b10000110100010011101001001011000000101000101011110;
        12'd38: TDATA = 50'b10000110100000011001000011011000000001000010000101;
        12'd39: TDATA = 50'b10000110011110010101001001010111111100111111001101;
        12'd40: TDATA = 50'b10000110011100010001001111010111111000111100011101;
        12'd41: TDATA = 50'b10000110011010001101011011010111110100111010000000;
        12'd42: TDATA = 50'b10000110011000001001101111010111110000110111111100;
        12'd43: TDATA = 50'b10000110010110000110000111010111101100110110000111;
        12'd44: TDATA = 50'b10000110010100000010100011010111101000110100011111;
        12'd45: TDATA = 50'b10000110010001111111001101010111100100110011011100;
        12'd46: TDATA = 50'b10000110001111111011111001010111100000110010101000;
        12'd47: TDATA = 50'b10000110001101111000101101010111011100110010000110;
        12'd48: TDATA = 50'b10000110001011110101011111010111011000110001101101;
        12'd49: TDATA = 50'b10000110001001110010100001010111010100110001111001;
        12'd50: TDATA = 50'b10000110000111101111100111010111010000110010010010;
        12'd51: TDATA = 50'b10000110000101101100101111010111001100110010111001;
        12'd52: TDATA = 50'b10000110000011101001111101010111001000110011110100;
        12'd53: TDATA = 50'b10000110000001100111010011010111000100110101001000;
        12'd54: TDATA = 50'b10000101111111100100110001010111000000110110101111;
        12'd55: TDATA = 50'b10000101111101100010010001010110111100111000100100;
        12'd56: TDATA = 50'b10000101111011011111111001010110111000111010110010;
        12'd57: TDATA = 50'b10000101111001011101100011010110110100111101001000;
        12'd58: TDATA = 50'b10000101110111011011010111010110110000111111111100;
        12'd59: TDATA = 50'b10000101110101011001001111010110101101000010111111;
        12'd60: TDATA = 50'b10000101110011010111010011010110101001000110100000;
        12'd61: TDATA = 50'b10000101110001010101010111010110100101001010001001;
        12'd62: TDATA = 50'b10000101101111010011100101010110100001001110001011;
        12'd63: TDATA = 50'b10000101101101010001110001010110011101010010010101;
        12'd64: TDATA = 50'b10000101101011010000001011010110011001010110111110;
        12'd65: TDATA = 50'b10000101101001001110101001010110010101011011111010;
        12'd66: TDATA = 50'b10000101100111001101001001010110010001100000111110;
        12'd67: TDATA = 50'b10000101100101001011110011010110001101100110100000;
        12'd68: TDATA = 50'b10000101100011001010100001010110001001101100010000;
        12'd69: TDATA = 50'b10000101100001001001010011010110000101110010001101;
        12'd70: TDATA = 50'b10000101011111001000001111010110000001111000101001;
        12'd71: TDATA = 50'b10000101011101000111001111010101111101111111010010;
        12'd72: TDATA = 50'b10000101011011000110011001010101111010000110010100;
        12'd73: TDATA = 50'b10000101011001000101100001010101110110001101011110;
        12'd74: TDATA = 50'b10000101010111000100110011010101110010010101000001;
        12'd75: TDATA = 50'b10000101010101000100001011010101101110011100110110;
        12'd76: TDATA = 50'b10000101010011000011100111010101101010100100111001;
        12'd77: TDATA = 50'b10000101010001000011001011010101100110101101010101;
        12'd78: TDATA = 50'b10000101001111000010110101010101100010110110000011;
        12'd79: TDATA = 50'b10000101001101000010100101010101011110111111000101;
        12'd80: TDATA = 50'b10000101001011000010010101010101011011001000001110;
        12'd81: TDATA = 50'b10000101001001000010010011010101010111010001111100;
        12'd82: TDATA = 50'b10000101000111000010001111010101010011011011101011;
        12'd83: TDATA = 50'b10000101000101000010010101010101001111100101110010;
        12'd84: TDATA = 50'b10000101000011000010100011010101001011110000010011;
        12'd85: TDATA = 50'b10000101000001000010110111010101000111111011000110;
        12'd86: TDATA = 50'b10000100111111000011001011010101000100000110000001;
        12'd87: TDATA = 50'b10000100111101000011101011010101000000010001011010;
        12'd88: TDATA = 50'b10000100111011000100001011010100111100011100111010;
        12'd89: TDATA = 50'b10000100111001000100110001010100111000101000101110;
        12'd90: TDATA = 50'b10000100110111000101011111010100110100110100111001;
        12'd91: TDATA = 50'b10000100110101000110010001010100110001000001010010;
        12'd92: TDATA = 50'b10000100110011000111001101010100101101001110000011;
        12'd93: TDATA = 50'b10000100110001001000001011010100101001011011000010;
        12'd94: TDATA = 50'b10000100101111001001010001010100100101101000011000;
        12'd95: TDATA = 50'b10000100101101001010011011010100100001110101111100;
        12'd96: TDATA = 50'b10000100101011001011101011010100011110000011110011;
        12'd97: TDATA = 50'b10000100101001001101000001010100011010010001111100;
        12'd98: TDATA = 50'b10000100100111001110100001010100010110100000011101;
        12'd99: TDATA = 50'b10000100100101001111111101010100010010101111000000;
        12'd100: TDATA = 50'b10000100100011010001100101010100001110111110000001;
        12'd101: TDATA = 50'b10000100100001010011001111010100001011001101001111;
        12'd102: TDATA = 50'b10000100011111010101000011010100000111011100110101;
        12'd103: TDATA = 50'b10000100011101010110111011010100000011101100101001;
        12'd104: TDATA = 50'b10000100011011011000110111010011111111111100101110;
        12'd105: TDATA = 50'b10000100011001011010110111010011111100001101000001;
        12'd106: TDATA = 50'b10000100010111011101000011010011111000011101110001;
        12'd107: TDATA = 50'b10000100010101011111010011010011110100101110101111;
        12'd108: TDATA = 50'b10000100010011100001100111010011110000111111111110;
        12'd109: TDATA = 50'b10000100010001100011111111010011101101010001011011;
        12'd110: TDATA = 50'b10000100001111100110011011010011101001100011000100;
        12'd111: TDATA = 50'b10000100001101101001000001010011100101110101001100;
        12'd112: TDATA = 50'b10000100001011101011101011010011100010000111011111;
        12'd113: TDATA = 50'b10000100001001101110011011010011011110011010000110;
        12'd114: TDATA = 50'b10000100000111110001010001010011011010101100111111;
        12'd115: TDATA = 50'b10000100000101110100001011010011010111000000000100;
        12'd116: TDATA = 50'b10000100000011110111001001010011010011010011011100;
        12'd117: TDATA = 50'b10000100000001111010010001010011001111100111001100;
        12'd118: TDATA = 50'b10000011111111111101011001010011001011111011000010;
        12'd119: TDATA = 50'b10000011111110000000110001010011001000001111011100;
        12'd120: TDATA = 50'b10000011111100000100000101010011000100100011111000;
        12'd121: TDATA = 50'b10000011111010000111011111010011000000111000100101;
        12'd122: TDATA = 50'b10000011111000001011000001010010111101001101101011;
        12'd123: TDATA = 50'b10000011110110001110100111010010111001100010111101;
        12'd124: TDATA = 50'b10000011110100010010010111010010110101111000100111;
        12'd125: TDATA = 50'b10000011110010010110000011010010110010001110010011;
        12'd126: TDATA = 50'b10000011110000011001111011010010101110100100011100;
        12'd127: TDATA = 50'b10000011101110011101111111010010101010111011000010;
        12'd128: TDATA = 50'b10000011101100100001111101010010100111010001100100;
        12'd129: TDATA = 50'b10000011101010100110000111010010100011101000100011;
        12'd130: TDATA = 50'b10000011101000101010010011010010011111111111101111;
        12'd131: TDATA = 50'b10000011100110101110100111010010011100010111001101;
        12'd132: TDATA = 50'b10000011100100110010111101010010011000101110110111;
        12'd133: TDATA = 50'b10000011100010110111011001010010010101000110110100;
        12'd134: TDATA = 50'b10000011100000111100000001010010010001011111001101;
        12'd135: TDATA = 50'b10000011011111000000101001010010001101110111101110;
        12'd136: TDATA = 50'b10000011011101000101010111010010001010010000100001;
        12'd137: TDATA = 50'b10000011011011001010000101010010000110101001011010;
        12'd138: TDATA = 50'b10000011011001001111000001010010000011000010110110;
        12'd139: TDATA = 50'b10000011010111010011111111010001111111011100011001;
        12'd140: TDATA = 50'b10000011010101011001000001010001111011110110001110;
        12'd141: TDATA = 50'b10000011010011011110010001010001111000010000100001;
        12'd142: TDATA = 50'b10000011010001100011011001010001110100101010101110;
        12'd143: TDATA = 50'b10000011001111101000101111010001110001000101011001;
        12'd144: TDATA = 50'b10000011001101101110000111010001101101100000010000;
        12'd145: TDATA = 50'b10000011001011110011100101010001101001111011011001;
        12'd146: TDATA = 50'b10000011001001111001001001010001100110010110110100;
        12'd147: TDATA = 50'b10000011000111111110101111010001100010110010011011;
        12'd148: TDATA = 50'b10000011000110000100011111010001011111001110011010;
        12'd149: TDATA = 50'b10000011000100001010001111010001011011101010011111;
        12'd150: TDATA = 50'b10000011000010010000001111010001011000000111000111;
        12'd151: TDATA = 50'b10000011000000010110000111010001010100100011101010;
        12'd152: TDATA = 50'b10000010111110011100001101010001010001000000101011;
        12'd153: TDATA = 50'b10000010111100100010010111010001001101011101111100;
        12'd154: TDATA = 50'b10000010111010101000101001010001001001111011100000;
        12'd155: TDATA = 50'b10000010111000101110111001010001000110011001001011;
        12'd156: TDATA = 50'b10000010110110110101010011010001000010110111001100;
        12'd157: TDATA = 50'b10000010110100111011110001010000111111010101011010;
        12'd158: TDATA = 50'b10000010110011000010010111010000111011110011111111;
        12'd159: TDATA = 50'b10000010110001001000111101010000111000010010101010;
        12'd160: TDATA = 50'b10000010101111001111101111010000110100110001110011;
        12'd161: TDATA = 50'b10000010101101010110011011010000110001010000110111;
        12'd162: TDATA = 50'b10000010101011011101011011010000101101110000101000;
        12'd163: TDATA = 50'b10000010101001100100010111010000101010010000010100;
        12'd164: TDATA = 50'b10000010100111101011010111010000100110110000010010;
        12'd165: TDATA = 50'b10000010100101110010100001010000100011010000101000;
        12'd166: TDATA = 50'b10000010100011111001101111010000011111110001001001;
        12'd167: TDATA = 50'b10000010100010000001000001010000011100010001111100;
        12'd168: TDATA = 50'b10000010100000001000011011010000011000110011000000;
        12'd169: TDATA = 50'b10000010011110001111111001010000010101010100010110;
        12'd170: TDATA = 50'b10000010011100010111011001010000010001110101110011;
        12'd171: TDATA = 50'b10000010011010011111000011010000001110010111101011;
        12'd172: TDATA = 50'b10000010011000100110110001010000001010111001110000;
        12'd173: TDATA = 50'b10000010010110101110100011010000000111011100000001;
        12'd174: TDATA = 50'b10000010010100110110011001010000000011111110100011;
        12'd175: TDATA = 50'b10000010010010111110010111010000000000100001010111;
        12'd176: TDATA = 50'b10000010010001000110011001001111111101000100011100;
        12'd177: TDATA = 50'b10000010001111001110011101001111111001100111100111;
        12'd178: TDATA = 50'b10000010001101010110101011001111110110001011001111;
        12'd179: TDATA = 50'b10000010001011011111000001001111110010101111001001;
        12'd180: TDATA = 50'b10000010001001100111010011001111101111010011000011;
        12'd181: TDATA = 50'b10000010000111101111110001001111101011110111011001;
        12'd182: TDATA = 50'b10000010000101111000001111001111101000011011110110;
        12'd183: TDATA = 50'b10000010000100000000110011001111100101000000100100;
        12'd184: TDATA = 50'b10000010000010001001011111001111100001100101101000;
        12'd185: TDATA = 50'b10000010000000010010001111001111011110001010111001;
        12'd186: TDATA = 50'b10000001111110011011000011001111011010110000010101;
        12'd187: TDATA = 50'b10000001111100100100000001001111010111010110001110;
        12'd188: TDATA = 50'b10000001111010101101000011001111010011111100010010;
        12'd189: TDATA = 50'b10000001111000110110001001001111010000100010100010;
        12'd190: TDATA = 50'b10000001110110111111010001001111001101001000111110;
        12'd191: TDATA = 50'b10000001110101001000011111001111001001101111101011;
        12'd192: TDATA = 50'b10000001110011010001110011001111000110010110101001;
        12'd193: TDATA = 50'b10000001110001011011001001001111000010111101110011;
        12'd194: TDATA = 50'b10000001101111100100100111001110111111100101001110;
        12'd195: TDATA = 50'b10000001101101101110001101001110111100001101000000;
        12'd196: TDATA = 50'b10000001101011110111110011001110111000110100111000;
        12'd197: TDATA = 50'b10000001101010000001100001001110110101011101000110;
        12'd198: TDATA = 50'b10000001101000001011010011001110110010000101100000;
        12'd199: TDATA = 50'b10000001100110010101001011001110101110101110001011;
        12'd200: TDATA = 50'b10000001100100011111000111001110101011010111000010;
        12'd201: TDATA = 50'b10000001100010101001000111001110101000000000001001;
        12'd202: TDATA = 50'b10000001100000110011001111001110100100101001100010;
        12'd203: TDATA = 50'b10000001011110111101011011001110100001010011001100;
        12'd204: TDATA = 50'b10000001011101000111101011001110011101111101000001;
        12'd205: TDATA = 50'b10000001011011010010000001001110011010100111001000;
        12'd206: TDATA = 50'b10000001011001011100011011001110010111010001011001;
        12'd207: TDATA = 50'b10000001010111100110111101001110010011111100000010;
        12'd208: TDATA = 50'b10000001010101110001100001001110010000100110110101;
        12'd209: TDATA = 50'b10000001010011111100001001001110001101010001110101;
        12'd210: TDATA = 50'b10000001010010000110110111001110001001111101000101;
        12'd211: TDATA = 50'b10000001010000010001101011001110000110101000100110;
        12'd212: TDATA = 50'b10000001001110011100100011001110000011010100010010;
        12'd213: TDATA = 50'b10000001001100100111011111001110000000000000010000;
        12'd214: TDATA = 50'b10000001001010110010100011001101111100101100011110;
        12'd215: TDATA = 50'b10000001001000111101101011001101111001011000111101;
        12'd216: TDATA = 50'b10000001000111001000110111001101110110000101101000;
        12'd217: TDATA = 50'b10000001000101010100001001001101110010110010100011;
        12'd218: TDATA = 50'b10000001000011011111011111001101101111011111101010;
        12'd219: TDATA = 50'b10000001000001101010111001001101101100001101000001;
        12'd220: TDATA = 50'b10000000111111110110011011001101101000111010101001;
        12'd221: TDATA = 50'b10000000111110000010000001001101100101101000100010;
        12'd222: TDATA = 50'b10000000111100001101101001001101100010010110100010;
        12'd223: TDATA = 50'b10000000111010011001011001001101011111000100110111;
        12'd224: TDATA = 50'b10000000111000100101001111001101011011110011011101;
        12'd225: TDATA = 50'b10000000110110110001000101001101011000100010001000;
        12'd226: TDATA = 50'b10000000110100111101000011001101010101010001001010;
        12'd227: TDATA = 50'b10000000110011001001001001001101010010000000011101;
        12'd228: TDATA = 50'b10000000110001010101010001001101001110101111111011;
        12'd229: TDATA = 50'b10000000101111100001011001001101001011011111011110;
        12'd230: TDATA = 50'b10000000101101101101101001001101001000001111011000;
        12'd231: TDATA = 50'b10000000101011111010000001001101000100111111100010;
        12'd232: TDATA = 50'b10000000101010000110011011001101000001101111111000;
        12'd233: TDATA = 50'b10000000101000010010111011001100111110100000011110;
        12'd234: TDATA = 50'b10000000100110011111100001001100111011010001010101;
        12'd235: TDATA = 50'b10000000100100101100001001001100111000000010010110;
        12'd236: TDATA = 50'b10000000100010111000111001001100110100110011101001;
        12'd237: TDATA = 50'b10000000100001000101101011001100110001100101000111;
        12'd238: TDATA = 50'b10000000011111010010100011001100101110010110110101;
        12'd239: TDATA = 50'b10000000011101011111100011001100101011001000111001;
        12'd240: TDATA = 50'b10000000011011101100100001001100100111111010111110;
        12'd241: TDATA = 50'b10000000011001111001101011001100100100101101011101;
        12'd242: TDATA = 50'b10000000011000000110110011001100100001011111111101;
        12'd243: TDATA = 50'b10000000010110010100000011001100011110010010110011;
        12'd244: TDATA = 50'b10000000010100100001011001001100011011000101111010;
        12'd245: TDATA = 50'b10000000010010101110110001001100010111111001001011;
        12'd246: TDATA = 50'b10000000010000111100010001001100010100101100101101;
        12'd247: TDATA = 50'b10000000001111001001110011001100010001100000011010;
        12'd248: TDATA = 50'b10000000001101010111011011001100001110010100010111;
        12'd249: TDATA = 50'b10000000001011100101001001001100001011001000100101;
        12'd250: TDATA = 50'b10000000001001110010111001001100000111111100111110;
        12'd251: TDATA = 50'b10000000001000000000110011001100000100110001101100;
        12'd252: TDATA = 50'b10000000000110001110101011001100000001100110011011;
        12'd253: TDATA = 50'b10000000000100011100110001001011111110011011101010;
        12'd254: TDATA = 50'b10000000000010101010110011001011111011010000111001;
        12'd255: TDATA = 50'b10000000000000111000111001001011111000000110010100;
        12'd256: TDATA = 50'b01111111111111000111001001001011110100111100000100;
        12'd257: TDATA = 50'b01111111111101010101011011001011110001110001111111;
        12'd258: TDATA = 50'b01111111111011100011110011001011101110101000001010;
        12'd259: TDATA = 50'b01111111111001110010010011001011101011011110101011;
        12'd260: TDATA = 50'b01111111111000000000110001001011101000010101001100;
        12'd261: TDATA = 50'b01111111110110001111011001001011100101001100000010;
        12'd262: TDATA = 50'b01111111110100011110000011001011100010000011000100;
        12'd263: TDATA = 50'b01111111110010101100101111001011011110111010010000;
        12'd264: TDATA = 50'b01111111110000111011100011001011011011110001101101;
        12'd265: TDATA = 50'b01111111101111001010011111001011011000101001011111;
        12'd266: TDATA = 50'b01111111101101011001010111001011010101100001010001;
        12'd267: TDATA = 50'b01111111101011101000011101001011010010011001011110;
        12'd268: TDATA = 50'b01111111101001110111100101001011001111010001110110;
        12'd269: TDATA = 50'b01111111101000000110101101001011001100001010010011;
        12'd270: TDATA = 50'b01111111100110010110000001001011001001000011001011;
        12'd271: TDATA = 50'b01111111100100100101010101001011000101111100001001;
        12'd272: TDATA = 50'b01111111100010110100101111001011000010110101010111;
        12'd273: TDATA = 50'b01111111100001000100001111001010111111101110110100;
        12'd274: TDATA = 50'b01111111011111010011101111001010111100101000011000;
        12'd275: TDATA = 50'b01111111011101100011010101001010111001100010001011;
        12'd276: TDATA = 50'b01111111011011110011000011001010110110011100010011;
        12'd277: TDATA = 50'b01111111011010000010110011001010110011010110100001;
        12'd278: TDATA = 50'b01111111011000010010100111001010110000010001000000;
        12'd279: TDATA = 50'b01111111010110100010011111001010101101001011101000;
        12'd280: TDATA = 50'b01111111010100110010100011001010101010000110101100;
        12'd281: TDATA = 50'b01111111010011000010100101001010100111000001101111;
        12'd282: TDATA = 50'b01111111010001010010101011001010100011111101000011;
        12'd283: TDATA = 50'b01111111001111100010111001001010100000111000100110;
        12'd284: TDATA = 50'b01111111001101110011001001001010011101110100010100;
        12'd285: TDATA = 50'b01111111001100000011011111001010011010110000010010;
        12'd286: TDATA = 50'b01111111001010010011110111001010010111101100011010;
        12'd287: TDATA = 50'b01111111001000100100010111001010010100101000110011;
        12'd288: TDATA = 50'b01111111000110110100111011001010010001100101011011;
        12'd289: TDATA = 50'b01111111000101000101100011001010001110100010001110;
        12'd290: TDATA = 50'b01111111000011010110001111001010001011011111001100;
        12'd291: TDATA = 50'b01111111000001100110111111001010001000011100011001;
        12'd292: TDATA = 50'b01111110111111110111110111001010000101011001110110;
        12'd293: TDATA = 50'b01111110111110001000110001001010000010010111011110;
        12'd294: TDATA = 50'b01111110111100011001110001001001111111010101010110;
        12'd295: TDATA = 50'b01111110111010101010110001001001111100010011010010;
        12'd296: TDATA = 50'b01111110111000111011111001001001111001010001100100;
        12'd297: TDATA = 50'b01111110110111001101000011001001110110001111111011;
        12'd298: TDATA = 50'b01111110110101011110010111001001110011001110101101;
        12'd299: TDATA = 50'b01111110110011101111101001001001110000001101011110;
        12'd300: TDATA = 50'b01111110110010000001000111001001101101001100101010;
        12'd301: TDATA = 50'b01111110110000010010100011001001101010001011110110;
        12'd302: TDATA = 50'b01111110101110100100001001001001100111001011011100;
        12'd303: TDATA = 50'b01111110101100110101110001001001100100001011000111;
        12'd304: TDATA = 50'b01111110101011000111011011001001100001001010111100;
        12'd305: TDATA = 50'b01111110101001011001001011001001011110001011000001;
        12'd306: TDATA = 50'b01111110100111101011000001001001011011001011010110;
        12'd307: TDATA = 50'b01111110100101111100111001001001011000001011110110;
        12'd308: TDATA = 50'b01111110100100001110111011001001010101001100101010;
        12'd309: TDATA = 50'b01111110100010100000110111001001010010001101011001;
        12'd310: TDATA = 50'b01111110100000110010111111001001001111001110100010;
        12'd311: TDATA = 50'b01111110011111000101010001001001001100001111111111;
        12'd312: TDATA = 50'b01111110011101010111011011001001001001010001011000;
        12'd313: TDATA = 50'b01111110011011101001101111001001000110010011000101;
        12'd314: TDATA = 50'b01111110011001111100001001001001000011010101000010;
        12'd315: TDATA = 50'b01111110011000001110100111001001000000010111001001;
        12'd316: TDATA = 50'b01111110010110100001001001001000111101011001100000;
        12'd317: TDATA = 50'b01111110010100110011101111001000111010011100000001;
        12'd318: TDATA = 50'b01111110010011000110011001001000110111011110101100;
        12'd319: TDATA = 50'b01111110010001011001000111001000110100100001100111;
        12'd320: TDATA = 50'b01111110001111101011111001001000110001100100101101;
        12'd321: TDATA = 50'b01111110001101111110110101001000101110101000000110;
        12'd322: TDATA = 50'b01111110001100010001101111001000101011101011100101;
        12'd323: TDATA = 50'b01111110001010100100110011001000101000101111011001;
        12'd324: TDATA = 50'b01111110001000110111110101001000100101110011001100;
        12'd325: TDATA = 50'b01111110000111001011000001001000100010110111011010;
        12'd326: TDATA = 50'b01111110000101011110001111001000011111111011101100;
        12'd327: TDATA = 50'b01111110000011110001011111001000011101000000001001;
        12'd328: TDATA = 50'b01111110000010000100110111001000011010000100111010;
        12'd329: TDATA = 50'b01111110000000011000010011001000010111001001110101;
        12'd330: TDATA = 50'b01111101111110101011101111001000010100001110110101;
        12'd331: TDATA = 50'b01111101111100111111010101001000010001010100001010;
        12'd332: TDATA = 50'b01111101111011010010111101001000001110011001101001;
        12'd333: TDATA = 50'b01111101111001100110100111001000001011011111010011;
        12'd334: TDATA = 50'b01111101110111111010011011001000001000100101010000;
        12'd335: TDATA = 50'b01111101110110001110001101001000000101101011001110;
        12'd336: TDATA = 50'b01111101110100100010001001001000000010110001100101;
        12'd337: TDATA = 50'b01111101110010110110000111000111111111111000000001;
        12'd338: TDATA = 50'b01111101110001001010001001000111111100111110101101;
        12'd339: TDATA = 50'b01111101101111011110001111000111111010000101100010;
        12'd340: TDATA = 50'b01111101101101110010011011000111110111001100100111;
        12'd341: TDATA = 50'b01111101101100000110101011000111110100010011110110;
        12'd342: TDATA = 50'b01111101101010011010111111000111110001011011010100;
        12'd343: TDATA = 50'b01111101101000101111010111000111101110100010111100;
        12'd344: TDATA = 50'b01111101100111000011101111000111101011101010101010;
        12'd345: TDATA = 50'b01111101100101011000010011000111101000110010110000;
        12'd346: TDATA = 50'b01111101100011101100110111000111100101111010111100;
        12'd347: TDATA = 50'b01111101100010000001100001000111100011000011010111;
        12'd348: TDATA = 50'b01111101100000010110001111000111100000001011111011;
        12'd349: TDATA = 50'b01111101011110101010111111000111011101010100101010;
        12'd350: TDATA = 50'b01111101011100111111110111000111011010011101101101;
        12'd351: TDATA = 50'b01111101011011010100110011000111010111100110111010;
        12'd352: TDATA = 50'b01111101011001101001101111000111010100110000001100;
        12'd353: TDATA = 50'b01111101010111111110110101000111010001111001110010;
        12'd354: TDATA = 50'b01111101010110010011111101000111001111000011100010;
        12'd355: TDATA = 50'b01111101010100101001000101000111001100001101010111;
        12'd356: TDATA = 50'b01111101010010111110011001000111001001010111100110;
        12'd357: TDATA = 50'b01111101010001010011101001000111000110100001110100;
        12'd358: TDATA = 50'b01111101001111101001000011000111000011101100010110;
        12'd359: TDATA = 50'b01111101001101111110100001000111000000110111000010;
        12'd360: TDATA = 50'b01111101001100010100000001000110111110000001111000;
        12'd361: TDATA = 50'b01111101001010101001100111000110111011001100111101;
        12'd362: TDATA = 50'b01111101001000111111001111000110111000011000001100;
        12'd363: TDATA = 50'b01111101000111010100111111000110110101100011101010;
        12'd364: TDATA = 50'b01111101000101101010101011000110110010101111000111;
        12'd365: TDATA = 50'b01111101000100000000100011000110101111111010111110;
        12'd366: TDATA = 50'b01111101000010010110011011000110101101000110111010;
        12'd367: TDATA = 50'b01111101000000101100011011000110101010010011001001;
        12'd368: TDATA = 50'b01111100111111000010011101000110100111011111011110;
        12'd369: TDATA = 50'b01111100111101011000100111000110100100101100000110;
        12'd370: TDATA = 50'b01111100111011101110110011000110100001111000111000;
        12'd371: TDATA = 50'b01111100111010000101000001000110011111000101101111;
        12'd372: TDATA = 50'b01111100111000011011010011000110011100010010110101;
        12'd373: TDATA = 50'b01111100110110110001101001000110011001100000000101;
        12'd374: TDATA = 50'b01111100110101001000001001000110010110101101101000;
        12'd375: TDATA = 50'b01111100110011011110100111000110010011111011010000;
        12'd376: TDATA = 50'b01111100110001110101001101000110010001001001000111;
        12'd377: TDATA = 50'b01111100110000001011110101000110001110010111001000;
        12'd378: TDATA = 50'b01111100101110100010011111000110001011100101010011;
        12'd379: TDATA = 50'b01111100101100111001010001000110001000110011101101;
        12'd380: TDATA = 50'b01111100101011010000000101000110000110000010010000;
        12'd381: TDATA = 50'b01111100101001100111000001000110000011010001000111;
        12'd382: TDATA = 50'b01111100100111111101111111000110000000100000000011;
        12'd383: TDATA = 50'b01111100100110010100111111000101111101101111001000;
        12'd384: TDATA = 50'b01111100100100101100000001000101111010111110010111;
        12'd385: TDATA = 50'b01111100100011000011001011000101111000001101110101;
        12'd386: TDATA = 50'b01111100100001011010011001000101110101011101100010;
        12'd387: TDATA = 50'b01111100011111110001101111000101110010101101011101;
        12'd388: TDATA = 50'b01111100011110001001000011000101101111111101011101;
        12'd389: TDATA = 50'b01111100011100100000011011000101101101001101100111;
        12'd390: TDATA = 50'b01111100011010110111111001000101101010011101111111;
        12'd391: TDATA = 50'b01111100011001001111011011000101100111101110100001;
        12'd392: TDATA = 50'b01111100010111100111000101000101100100111111010111;
        12'd393: TDATA = 50'b01111100010101111110101111000101100010010000010001;
        12'd394: TDATA = 50'b01111100010100010110011111000101011111100001011010;
        12'd395: TDATA = 50'b01111100010010101110001111000101011100110010101000;
        12'd396: TDATA = 50'b01111100010001000110000111000101011010000100001001;
        12'd397: TDATA = 50'b01111100001111011110000011000101010111010101110100;
        12'd398: TDATA = 50'b01111100001101110101111111000101010100100111100011;
        12'd399: TDATA = 50'b01111100001100001110000101000101010001111001100110;
        12'd400: TDATA = 50'b01111100001010100110001101000101001111001011110011;
        12'd401: TDATA = 50'b01111100001000111110010101000101001100011110000100;
        12'd402: TDATA = 50'b01111100000111010110101001000101001001110000101101;
        12'd403: TDATA = 50'b01111100000101101110111001000101000111000011010110;
        12'd404: TDATA = 50'b01111100000100000111010001000101000100010110001110;
        12'd405: TDATA = 50'b01111100000010011111101011000101000001101001001111;
        12'd406: TDATA = 50'b01111100000000111000001011000100111110111100011111;
        12'd407: TDATA = 50'b01111011111111010000110001000100111100001111111110;
        12'd408: TDATA = 50'b01111011111101101001010111000100111001100011100000;
        12'd409: TDATA = 50'b01111011111100000010000011000100110110110111010010;
        12'd410: TDATA = 50'b01111011111010011010110001000100110100001011001100;
        12'd411: TDATA = 50'b01111011111000110011100111000100110001011111010110;
        12'd412: TDATA = 50'b01111011110111001100011111000100101110110011101001;
        12'd413: TDATA = 50'b01111011110101100101011001000100101100001000000101;
        12'd414: TDATA = 50'b01111011110011111110010111000100101001011100101010;
        12'd415: TDATA = 50'b01111011110010010111011011000100100110110001011110;
        12'd416: TDATA = 50'b01111011110000110000100011000100100100000110011100;
        12'd417: TDATA = 50'b01111011101111001001101111000100100001011011101000;
        12'd418: TDATA = 50'b01111011101101100010111111000100011110110000111101;
        12'd419: TDATA = 50'b01111011101011111100010011000100011100000110011100;
        12'd420: TDATA = 50'b01111011101010010101101111000100011001011100001110;
        12'd421: TDATA = 50'b01111011101000101111000111000100010110110010000000;
        12'd422: TDATA = 50'b01111011100111001000100111000100010100001000000000;
        12'd423: TDATA = 50'b01111011100101100010001011000100010001011110001110;
        12'd424: TDATA = 50'b01111011100011111011110011000100001110110100100101;
        12'd425: TDATA = 50'b01111011100010010101011111000100001100001011000110;
        12'd426: TDATA = 50'b01111011100000101111001101000100001001100001110001;
        12'd427: TDATA = 50'b01111011011111001001000011000100000110111000101110;
        12'd428: TDATA = 50'b01111011011101100010111011000100000100001111110000;
        12'd429: TDATA = 50'b01111011011011111100110101000100000001100110111011;
        12'd430: TDATA = 50'b01111011011010010110110101000011111110111110010101;
        12'd431: TDATA = 50'b01111011011000110000110111000011111100010101111000;
        12'd432: TDATA = 50'b01111011010111001011000001000011111001101101101001;
        12'd433: TDATA = 50'b01111011010101100101001001000011110111000101011110;
        12'd434: TDATA = 50'b01111011010011111111011011000011110100011101100111;
        12'd435: TDATA = 50'b01111011010010011001101011000011110001110101101111;
        12'd436: TDATA = 50'b01111011010000110100000011000011101111001110001011;
        12'd437: TDATA = 50'b01111011001111001110100011000011101100100110111001;
        12'd438: TDATA = 50'b01111011001101101000111111000011101001111111100010;
        12'd439: TDATA = 50'b01111011001100000011011111000011100111011000011001;
        12'd440: TDATA = 50'b01111011001010011110001001000011100100110001100011;
        12'd441: TDATA = 50'b01111011001000111000110011000011100010001010110001;
        12'd442: TDATA = 50'b01111011000111010011100011000011011111100100001101;
        12'd443: TDATA = 50'b01111011000101101110010111000011011100111101110011;
        12'd444: TDATA = 50'b01111011000100001001001001000011011010010111011101;
        12'd445: TDATA = 50'b01111011000010100100001001000011010111110001011111;
        12'd446: TDATA = 50'b01111011000000111111000101000011010101001011100001;
        12'd447: TDATA = 50'b01111010111111011010000111000011010010100101110000;
        12'd448: TDATA = 50'b01111010111101110101001011000011010000000000001001;
        12'd449: TDATA = 50'b01111010111100010000010111000011001101011010101111;
        12'd450: TDATA = 50'b01111010111010101011100101000011001010110101011111;
        12'd451: TDATA = 50'b01111010111001000110111001000011001000010000011101;
        12'd452: TDATA = 50'b01111010110111100010001101000011000101101011011111;
        12'd453: TDATA = 50'b01111010110101111101100111000011000011000110101111;
        12'd454: TDATA = 50'b01111010110100011001000011000011000000100010001001;
        12'd455: TDATA = 50'b01111010110010110100100111000010111101111101110000;
        12'd456: TDATA = 50'b01111010110001010000001001000010111011011001011100;
        12'd457: TDATA = 50'b01111010101111101011101111000010111000110101010000;
        12'd458: TDATA = 50'b01111010101110000111011111000010110110010001011000;
        12'd459: TDATA = 50'b01111010101100100011001011000010110011101101011111;
        12'd460: TDATA = 50'b01111010101010111111000011000010110001001001111101;
        12'd461: TDATA = 50'b01111010101001011010110111000010101110100110011011;
        12'd462: TDATA = 50'b01111010100111110110111001000010101100000011010001;
        12'd463: TDATA = 50'b01111010100110010010110111000010101001100000000110;
        12'd464: TDATA = 50'b01111010100100101110111011000010100110111101001001;
        12'd465: TDATA = 50'b01111010100011001011000001000010100100011010010101;
        12'd466: TDATA = 50'b01111010100001100111001111000010100001110111101110;
        12'd467: TDATA = 50'b01111010100000000011011111000010011111010101010001;
        12'd468: TDATA = 50'b01111010011110011111101111000010011100110010111000;
        12'd469: TDATA = 50'b01111010011100111100000111000010011010010000110010;
        12'd470: TDATA = 50'b01111010011011011000100011000010010111101110110101;
        12'd471: TDATA = 50'b01111010011001110100111111000010010101001100111100;
        12'd472: TDATA = 50'b01111010011000010001100001000010010010101011010000;
        12'd473: TDATA = 50'b01111010010110101110001001000010010000001001110011;
        12'd474: TDATA = 50'b01111010010101001010110001000010001101101000011010;
        12'd475: TDATA = 50'b01111010010011100111011101000010001011000111001001;
        12'd476: TDATA = 50'b01111010010010000100010001000010001000100110001100;
        12'd477: TDATA = 50'b01111010010000100001000101000010000110000101010010;
        12'd478: TDATA = 50'b01111010001110111101111111000010000011100100100110;
        12'd479: TDATA = 50'b01111010001101011010111011000010000001000100000011;
        12'd480: TDATA = 50'b01111010001011110111111001000001111110100011100101;
        12'd481: TDATA = 50'b01111010001010010100111111000001111100000011011000;
        12'd482: TDATA = 50'b01111010001000110010000101000001111001100011010000;
        12'd483: TDATA = 50'b01111010000111001111010001000001110111000011010110;
        12'd484: TDATA = 50'b01111010000101101100011111000001110100100011100100;
        12'd485: TDATA = 50'b01111010000100001001110001000001110010000011111100;
        12'd486: TDATA = 50'b01111010000010100111001001000001101111100100100001;
        12'd487: TDATA = 50'b01111010000001000100100101000001101101000101001111;
        12'd488: TDATA = 50'b01111001111111100001111111000001101010100110000001;
        12'd489: TDATA = 50'b01111001111101111111100011000001101000000111000110;
        12'd490: TDATA = 50'b01111001111100011101001011000001100101101000010011;
        12'd491: TDATA = 50'b01111001111010111010110101000001100011001001101010;
        12'd492: TDATA = 50'b01111001111001011000100001000001100000101011001001;
        12'd493: TDATA = 50'b01111001110111110110010001000001011110001100110001;
        12'd494: TDATA = 50'b01111001110110010100000111000001011011101110100110;
        12'd495: TDATA = 50'b01111001110100110010000001000001011001010000100101;
        12'd496: TDATA = 50'b01111001110011001111111101000001010110110010101100;
        12'd497: TDATA = 50'b01111001110001101101111011000001010100010100111100;
        12'd498: TDATA = 50'b01111001110000001100000001000001010001110111011010;
        12'd499: TDATA = 50'b01111001101110101010000011000001001111011001110111;
        12'd500: TDATA = 50'b01111001101101001000010001000001001100111100101011;
        12'd501: TDATA = 50'b01111001101011100110011111000001001010011111100011;
        12'd502: TDATA = 50'b01111001101010000100101111000001001000000010100011;
        12'd503: TDATA = 50'b01111001101000100011001001000001000101100101110110;
        12'd504: TDATA = 50'b01111001100111000001100001000001000011001001001001;
        12'd505: TDATA = 50'b01111001100101011111111011000001000000101100100100;
        12'd506: TDATA = 50'b01111001100011111110100001000000111110010000010110;
        12'd507: TDATA = 50'b01111001100010011101000001000000111011110100000010;
        12'd508: TDATA = 50'b01111001100000111011101001000000111001011000000001;
        12'd509: TDATA = 50'b01111001011111011010010011000000110110111100000100;
        12'd510: TDATA = 50'b01111001011101111001000101000000110100100000011001;
        12'd511: TDATA = 50'b01111001011100010111110111000000110010000100110010;
        12'd512: TDATA = 50'b01111001011010110110101111000000101111101001011000;
        12'd513: TDATA = 50'b01111001011001010101101001000000101101001110000111;
        12'd514: TDATA = 50'b01111001010111110100100111000000101010110010111111;
        12'd515: TDATA = 50'b01111001010110010011101011000000101000011000000100;
        12'd516: TDATA = 50'b01111001010100110010101101000000100101111101001001;
        12'd517: TDATA = 50'b01111001010011010001111001000000100011100010100100;
        12'd518: TDATA = 50'b01111001010001110001000011000000100001000111111110;
        12'd519: TDATA = 50'b01111001010000010000010111000000011110101101101011;
        12'd520: TDATA = 50'b01111001001110101111100111000000011100010011010111;
        12'd521: TDATA = 50'b01111001001101001110111111000000011001111001010100;
        12'd522: TDATA = 50'b01111001001011101110011011000000010111011111011011;
        12'd523: TDATA = 50'b01111001001010001101110111000000010101000101100101;
        12'd524: TDATA = 50'b01111001001000101101011001000000010010101011111101;
        12'd525: TDATA = 50'b01111001000111001101000001000000010000010010100010;
        12'd526: TDATA = 50'b01111001000101101100101001000000001101111001001011;
        12'd527: TDATA = 50'b01111001000100001100010101000000001011011111111100;
        12'd528: TDATA = 50'b01111001000010101100001001000000001001000111000000;
        12'd529: TDATA = 50'b01111001000001001011111001000000000110101110000010;
        12'd530: TDATA = 50'b01111000111111101011110011000000000100010101010111;
        12'd531: TDATA = 50'b01111000111110001011110001000000000001111100110100;
        12'd532: TDATA = 50'b01111000111100101011101010111111111111100100010001;
        12'd533: TDATA = 50'b01111000111011001011110000111111111101001100000100;
        12'd534: TDATA = 50'b01111000111001101011110110111111111010110011111011;
        12'd535: TDATA = 50'b01111000111000001011111110111111111000011011111010;
        12'd536: TDATA = 50'b01111000110110101100001110111111110110000100000111;
        12'd537: TDATA = 50'b01111000110101001100011010111111110011101100010010;
        12'd538: TDATA = 50'b01111000110011101100101110111111110001010100110000;
        12'd539: TDATA = 50'b01111000110010001101000110111111101110111101010110;
        12'd540: TDATA = 50'b01111000110000101101100010111111101100100110000101;
        12'd541: TDATA = 50'b01111000101111001110000010111111101010001111000001;
        12'd542: TDATA = 50'b01111000101101101110100100111111100111111000000001;
        12'd543: TDATA = 50'b01111000101100001111001010111111100101100001001101;
        12'd544: TDATA = 50'b01111000101010101111110010111111100011001010011110;
        12'd545: TDATA = 50'b01111000101001010000100010111111100000110100000001;
        12'd546: TDATA = 50'b01111000100111110001010010111111011110011101100111;
        12'd547: TDATA = 50'b01111000100110010010001000111111011100000111011010;
        12'd548: TDATA = 50'b01111000100100110010111110111111011001110001010001;
        12'd549: TDATA = 50'b01111000100011010011110110111111010111011011010001;
        12'd550: TDATA = 50'b01111000100001110100110110111111010101000101011110;
        12'd551: TDATA = 50'b01111000100000010101111010111111010010101111110111;
        12'd552: TDATA = 50'b01111000011110110111000000111111010000011010010101;
        12'd553: TDATA = 50'b01111000011101011000001000111111001110000100111011;
        12'd554: TDATA = 50'b01111000011011111001010110111111001011101111101110;
        12'd555: TDATA = 50'b01111000011010011010100100111111001001011010100101;
        12'd556: TDATA = 50'b01111000011000111011111000111111000111000101101001;
        12'd557: TDATA = 50'b01111000010111011101001110111111000100110000110101;
        12'd558: TDATA = 50'b01111000010101111110101000111111000010011100001001;
        12'd559: TDATA = 50'b01111000010100100000001000111111000000000111101011;
        12'd560: TDATA = 50'b01111000010011000001101000111110111101110011010000;
        12'd561: TDATA = 50'b01111000010001100011001110111110111011011111000011;
        12'd562: TDATA = 50'b01111000010000000100111000111110111001001010111101;
        12'd563: TDATA = 50'b01111000001110100110100000111110110110110110111100;
        12'd564: TDATA = 50'b01111000001101001000010110111110110100100011010000;
        12'd565: TDATA = 50'b01111000001011101010000010111110110010001111011011;
        12'd566: TDATA = 50'b01111000001010001011111010111110101111111011111011;
        12'd567: TDATA = 50'b01111000001000101101111000111110101101101000101001;
        12'd568: TDATA = 50'b01111000000111001111110010111110101011010101010110;
        12'd569: TDATA = 50'b01111000000101110001110100111110101001000010001111;
        12'd570: TDATA = 50'b01111000000100010011111010111110100110101111010110;
        12'd571: TDATA = 50'b01111000000010110101111110111110100100011100011100;
        12'd572: TDATA = 50'b01111000000001011000001100111110100010001001110011;
        12'd573: TDATA = 50'b01110111111111111010011000111110011111110111001110;
        12'd574: TDATA = 50'b01110111111110011100101000111110011101100100110000;
        12'd575: TDATA = 50'b01110111111100111110111110111110011011010010100000;
        12'd576: TDATA = 50'b01110111111011100001011010111110011001000000011101;
        12'd577: TDATA = 50'b01110111111010000011110100111110010110101110011001;
        12'd578: TDATA = 50'b01110111111000100110010110111110010100011100100110;
        12'd579: TDATA = 50'b01110111110111001000111010111110010010001010111100;
        12'd580: TDATA = 50'b01110111110101101011100000111110001111111001010101;
        12'd581: TDATA = 50'b01110111110100001110001000111110001101100111110110;
        12'd582: TDATA = 50'b01110111110010110000110110111110001011010110100101;
        12'd583: TDATA = 50'b01110111110001010011100100111110001001000101010110;
        12'd584: TDATA = 50'b01110111101111110110011010111110000110110100011010;
        12'd585: TDATA = 50'b01110111101110011001010010111110000100100011100001;
        12'd586: TDATA = 50'b01110111101100111100001100111110000010010010110000;
        12'd587: TDATA = 50'b01110111101011011111001100111110000000000010001100;
        12'd588: TDATA = 50'b01110111101010000010001100111101111101110001101011;
        12'd589: TDATA = 50'b01110111101000100101001110111101111011100001010010;
        12'd590: TDATA = 50'b01110111100111001000011010111101111001010001001011;
        12'd591: TDATA = 50'b01110111100101101011100110111101110111000001001000;
        12'd592: TDATA = 50'b01110111100100001110110110111101110100110001001100;
        12'd593: TDATA = 50'b01110111100010110010001000111101110010100001011001;
        12'd594: TDATA = 50'b01110111100001010101100000111101110000010001110011;
        12'd595: TDATA = 50'b01110111011111111000111000111101101110000010010000;
        12'd596: TDATA = 50'b01110111011110011100010010111101101011110010110101;
        12'd597: TDATA = 50'b01110111011100111111110100111101101001100011100111;
        12'd598: TDATA = 50'b01110111011011100011011000111101100111010100100001;
        12'd599: TDATA = 50'b01110111011010000110111100111101100101000101011111;
        12'd600: TDATA = 50'b01110111011000101010101000111101100010110110101110;
        12'd601: TDATA = 50'b01110111010111001110010110111101100000101000000000;
        12'd602: TDATA = 50'b01110111010101110010000110111101011110011001011010;
        12'd603: TDATA = 50'b01110111010100010101111000111101011100001010111101;
        12'd604: TDATA = 50'b01110111010010111001101110111101011001111100100111;
        12'd605: TDATA = 50'b01110111010001011101101110111101010111101110100011;
        12'd606: TDATA = 50'b01110111010000000001100110111101010101100000011001;
        12'd607: TDATA = 50'b01110111001110100101101100111101010011010010100101;
        12'd608: TDATA = 50'b01110111001101001001110000111101010001000100110101;
        12'd609: TDATA = 50'b01110111001011101101111000111101001110110111001100;
        12'd610: TDATA = 50'b01110111001010010010000100111101001100101001101100;
        12'd611: TDATA = 50'b01110111001000110110010010111101001010011100010011;
        12'd612: TDATA = 50'b01110111000111011010100010111101001000001111000011;
        12'd613: TDATA = 50'b01110111000101111110111010111101000110000001111111;
        12'd614: TDATA = 50'b01110111000100100011010000111101000011110100111111;
        12'd615: TDATA = 50'b01110111000011000111101110111101000001101000001011;
        12'd616: TDATA = 50'b01110111000001101100001110111100111111011011011111;
        12'd617: TDATA = 50'b01110111000000010000110000111100111101001110111011;
        12'd618: TDATA = 50'b01110110111110110101010100111100111011000010011011;
        12'd619: TDATA = 50'b01110110111101011010000000111100111000110110001011;
        12'd620: TDATA = 50'b01110110111011111110101000111100110110101001111011;
        12'd621: TDATA = 50'b01110110111010100011011110111100110100011110000000;
        12'd622: TDATA = 50'b01110110111001001000001010111100110010010001111011;
        12'd623: TDATA = 50'b01110110110111101101000010111100110000000110001100;
        12'd624: TDATA = 50'b01110110110110010001111010111100101101111010011111;
        12'd625: TDATA = 50'b01110110110100110110111010111100101011101111000100;
        12'd626: TDATA = 50'b01110110110011011011111000111100101001100011101000;
        12'd627: TDATA = 50'b01110110110010000001000000111100100111011000011101;
        12'd628: TDATA = 50'b01110110110000100110000100111100100101001101010001;
        12'd629: TDATA = 50'b01110110101111001011001110111100100011000010010001;
        12'd630: TDATA = 50'b01110110101101110000011010111100100000110111011001;
        12'd631: TDATA = 50'b01110110101100010101101110111100011110101100101110;
        12'd632: TDATA = 50'b01110110101010111010111110111100011100100010000001;
        12'd633: TDATA = 50'b01110110101001100000010110111100011010010111100101;
        12'd634: TDATA = 50'b01110110101000000101110000111100011000001101001101;
        12'd635: TDATA = 50'b01110110100110101011001100111100010110000010111100;
        12'd636: TDATA = 50'b01110110100101010000101110111100010011111000111001;
        12'd637: TDATA = 50'b01110110100011110110010010111100010001101110111100;
        12'd638: TDATA = 50'b01110110100010011011111000111100001111100101000100;
        12'd639: TDATA = 50'b01110110100001000001100010111100001101011011010111;
        12'd640: TDATA = 50'b01110110011111100111010000111100001011010001110011;
        12'd641: TDATA = 50'b01110110011110001100111110111100001001001000010001;
        12'd642: TDATA = 50'b01110110011100110010110110111100000110111111000001;
        12'd643: TDATA = 50'b01110110011011011000101010111100000100110101101111;
        12'd644: TDATA = 50'b01110110011001111110100100111100000010101100101010;
        12'd645: TDATA = 50'b01110110011000100100100100111100000000100011110001;
        12'd646: TDATA = 50'b01110110010111001010100100111011111110011010111100;
        12'd647: TDATA = 50'b01110110010101110000100110111011111100010010001110;
        12'd648: TDATA = 50'b01110110010100010110110000111011111010001001101100;
        12'd649: TDATA = 50'b01110110010010111100111000111011111000000001001110;
        12'd650: TDATA = 50'b01110110010001100011001000111011110101111000111100;
        12'd651: TDATA = 50'b01110110010000001001010110111011110011110000101110;
        12'd652: TDATA = 50'b01110110001110101111101100111011110001101000101100;
        12'd653: TDATA = 50'b01110110001101010110000000111011101111100000101100;
        12'd654: TDATA = 50'b01110110001011111100011110111011101101011000111110;
        12'd655: TDATA = 50'b01110110001010100010110110111011101011010001001010;
        12'd656: TDATA = 50'b01110110001001001001011010111011101001001001101011;
        12'd657: TDATA = 50'b01110110000111101111111110111011100111000010010000;
        12'd658: TDATA = 50'b01110110000110010110101000111011100100111011000001;
        12'd659: TDATA = 50'b01110110000100111101010010111011100010110011110101;
        12'd660: TDATA = 50'b01110110000011100100000000111011100000101100110001;
        12'd661: TDATA = 50'b01110110000010001010110000111011011110100101110100;
        12'd662: TDATA = 50'b01110110000000110001100010111011011100011110111111;
        12'd663: TDATA = 50'b01110101111111011000011000111011011010011000010010;
        12'd664: TDATA = 50'b01110101111101111111001110111011011000010001101000;
        12'd665: TDATA = 50'b01110101111100100110010000111011010110001011010100;
        12'd666: TDATA = 50'b01110101111011001101010010111011010100000101000010;
        12'd667: TDATA = 50'b01110101111001110100010010111011010001111110101111;
        12'd668: TDATA = 50'b01110101111000011011011010111011001111111000101101;
        12'd669: TDATA = 50'b01110101110111000010101000111011001101110010111000;
        12'd670: TDATA = 50'b01110101110101101001110000111011001011101100111100;
        12'd671: TDATA = 50'b01110101110100010001000000111011001001100111010001;
        12'd672: TDATA = 50'b01110101110010111000010010111011000111100001101001;
        12'd673: TDATA = 50'b01110101110001011111101000111011000101011100001101;
        12'd674: TDATA = 50'b01110101110000000111000110111011000011010110111101;
        12'd675: TDATA = 50'b01110101101110101110100010111011000001010001110001;
        12'd676: TDATA = 50'b01110101101101010110000000111010111111001100101000;
        12'd677: TDATA = 50'b01110101101011111101100110111010111101000111101111;
        12'd678: TDATA = 50'b01110101101010100101001000111010111011000010110101;
        12'd679: TDATA = 50'b01110101101001001100110010111010111000111110000111;
        12'd680: TDATA = 50'b01110101100111110100011110111010110110111001100001;
        12'd681: TDATA = 50'b01110101100110011100001010111010110100110100111110;
        12'd682: TDATA = 50'b01110101100101000011111110111010110010110000101011;
        12'd683: TDATA = 50'b01110101100011101011110110111010110000101100100000;
        12'd684: TDATA = 50'b01110101100010010011101110111010101110101000011000;
        12'd685: TDATA = 50'b01110101100000111011100110111010101100100100010011;
        12'd686: TDATA = 50'b01110101011111100011101010111010101010100000100100;
        12'd687: TDATA = 50'b01110101011110001011101000111010101000011100101110;
        12'd688: TDATA = 50'b01110101011100110011110000111010100110011001001001;
        12'd689: TDATA = 50'b01110101011011011011110100111010100100010101100011;
        12'd690: TDATA = 50'b01110101011010000100000000111010100010010010001101;
        12'd691: TDATA = 50'b01110101011000101100010000111010100000001110111110;
        12'd692: TDATA = 50'b01110101010111010100100000111010011110001011110011;
        12'd693: TDATA = 50'b01110101010101111100110100111010011100001000101111;
        12'd694: TDATA = 50'b01110101010100100101001010111010011010000101110011;
        12'd695: TDATA = 50'b01110101010011001101100110111010011000000011000011;
        12'd696: TDATA = 50'b01110101010001110110000010111010010110000000010110;
        12'd697: TDATA = 50'b01110101010000011110100100111010010011111101110101;
        12'd698: TDATA = 50'b01110101001111000111001000111010010001111011011011;
        12'd699: TDATA = 50'b01110101001101101111110000111010001111111001001001;
        12'd700: TDATA = 50'b01110101001100011000011000111010001101110110111010;
        12'd701: TDATA = 50'b01110101001011000001000100111010001011110100110010;
        12'd702: TDATA = 50'b01110101001001101001111000111010001001110010111011;
        12'd703: TDATA = 50'b01110101001000010010101000111010000111110001000010;
        12'd704: TDATA = 50'b01110101000110111011100000111010000101101111010110;
        12'd705: TDATA = 50'b01110101000101100100010100111010000011101101101000;
        12'd706: TDATA = 50'b01110101000100001101010100111010000001101100001110;
        12'd707: TDATA = 50'b01110101000010110110010000111001111111101010110100;
        12'd708: TDATA = 50'b01110101000001011111010100111001111101101001100101;
        12'd709: TDATA = 50'b01110101000000001000010110111001111011101000011001;
        12'd710: TDATA = 50'b01110100111110110001100000111001111001100111011001;
        12'd711: TDATA = 50'b01110100111101011010101100111001110111100110100001;
        12'd712: TDATA = 50'b01110100111100000011111010111001110101100101110000;
        12'd713: TDATA = 50'b01110100111010101101001010111001110011100101000010;
        12'd714: TDATA = 50'b01110100111001010110011110111001110001100100100000;
        12'd715: TDATA = 50'b01110100110111111111110110111001101111100100000101;
        12'd716: TDATA = 50'b01110100110110101001001110111001101101100011101101;
        12'd717: TDATA = 50'b01110100110101010010110000111001101011100011100110;
        12'd718: TDATA = 50'b01110100110011111100001110111001101001100011011101;
        12'd719: TDATA = 50'b01110100110010100101101110111001100111100011011100;
        12'd720: TDATA = 50'b01110100110001001111011000111001100101100011101010;
        12'd721: TDATA = 50'b01110100101111111001000010111001100011100011111100;
        12'd722: TDATA = 50'b01110100101110100010101010111001100001100100001100;
        12'd723: TDATA = 50'b01110100101101001100011010111001011111100100101101;
        12'd724: TDATA = 50'b01110100101011110110010000111001011101100101011001;
        12'd725: TDATA = 50'b01110100101010100000000010111001011011100110000100;
        12'd726: TDATA = 50'b01110100101001001001111000111001011001100110110110;
        12'd727: TDATA = 50'b01110100100111110011111000111001010111100111111001;
        12'd728: TDATA = 50'b01110100100110011101110100111001010101101000111010;
        12'd729: TDATA = 50'b01110100100101000111110110111001010011101010000110;
        12'd730: TDATA = 50'b01110100100011110001111010111001010001101011011010;
        12'd731: TDATA = 50'b01110100100010011100000010111001001111101100110110;
        12'd732: TDATA = 50'b01110100100001000110001010111001001101101110010100;
        12'd733: TDATA = 50'b01110100011111110000010110111001001011101111111010;
        12'd734: TDATA = 50'b01110100011110011010100110111001001001110001101011;
        12'd735: TDATA = 50'b01110100011101000100111010111001000111110011100100;
        12'd736: TDATA = 50'b01110100011011101111001110111001000101110101011111;
        12'd737: TDATA = 50'b01110100011010011001101000111001000011110111100111;
        12'd738: TDATA = 50'b01110100011001000100000110111001000001111001110101;
        12'd739: TDATA = 50'b01110100010111101110100010111000111111111100000111;
        12'd740: TDATA = 50'b01110100010110011001000110111000111101111110100100;
        12'd741: TDATA = 50'b01110100010101000011101000111000111100000001000100;
        12'd742: TDATA = 50'b01110100010011101110001110111000111010000011101011;
        12'd743: TDATA = 50'b01110100010010011000111010111000111000000110011110;
        12'd744: TDATA = 50'b01110100010001000011100110111000110110001001010100;
        12'd745: TDATA = 50'b01110100001111101110010110111000110100001100010001;
        12'd746: TDATA = 50'b01110100001110011001001110111000110010001111011111;
        12'd747: TDATA = 50'b01110100001101000100000010111000110000010010101010;
        12'd748: TDATA = 50'b01110100001011101110111010111000101110010101111101;
        12'd749: TDATA = 50'b01110100001010011001110110111000101100011001011000;
        12'd750: TDATA = 50'b01110100001001000100110100111000101010011100111001;
        12'd751: TDATA = 50'b01110100000111101111111010111000101000100000101011;
        12'd752: TDATA = 50'b01110100000110011010111100111000100110100100010110;
        12'd753: TDATA = 50'b01110100000101000110000010111000100100101000001101;
        12'd754: TDATA = 50'b01110100000011110001010000111000100010101100010000;
        12'd755: TDATA = 50'b01110100000010011100011010111000100000110000010001;
        12'd756: TDATA = 50'b01110100000001000111101010111000011110110100011110;
        12'd757: TDATA = 50'b01110011111111110011000000111000011100111000110110;
        12'd758: TDATA = 50'b01110011111110011110010110111000011010111101010001;
        12'd759: TDATA = 50'b01110011111101001001101110111000011001000001110100;
        12'd760: TDATA = 50'b01110011111011110101001010111000010111000110011101;
        12'd761: TDATA = 50'b01110011111010100000100110111000010101001011001010;
        12'd762: TDATA = 50'b01110011111001001100001000111000010011010000000010;
        12'd763: TDATA = 50'b01110011110111110111110000111000010001010101000101;
        12'd764: TDATA = 50'b01110011110110100011010110111000001111011010000111;
        12'd765: TDATA = 50'b01110011110101001111000000111000001101011111010101;
        12'd766: TDATA = 50'b01110011110011111010101100111000001011100100100101;
        12'd767: TDATA = 50'b01110011110010100110100000111000001001101010000101;
        12'd768: TDATA = 50'b01110011110001010010010000111000000111101111100011;
        12'd769: TDATA = 50'b01110011101111111110001000111000000101110101001101;
        12'd770: TDATA = 50'b01110011101110101001111110111000000011111010111010;
        12'd771: TDATA = 50'b01110011101101010101111100111000000010000000110011;
        12'd772: TDATA = 50'b01110011101100000001111000111000000000000110101110;
        12'd773: TDATA = 50'b01110011101010101101111000110111111110001100110000;
        12'd774: TDATA = 50'b01110011101001011001111110110111111100010010111110;
        12'd775: TDATA = 50'b01110011101000000110001000110111111010011001010010;
        12'd776: TDATA = 50'b01110011100110110010001110110111111000011111100110;
        12'd777: TDATA = 50'b01110011100101011110011010110111110110100110000100;
        12'd778: TDATA = 50'b01110011100100001010101100110111110100101100101111;
        12'd779: TDATA = 50'b01110011100010110110111110110111110010110011011011;
        12'd780: TDATA = 50'b01110011100001100011010110110111110000111010010100;
        12'd781: TDATA = 50'b01110011100000001111101010110111101111000001001010;
        12'd782: TDATA = 50'b01110011011110111100000110110111101101001000001100;
        12'd783: TDATA = 50'b01110011011101101000100100110111101011001111010110;
        12'd784: TDATA = 50'b01110011011100010101000010110111101001010110100010;
        12'd785: TDATA = 50'b01110011011011000001101000110111100111011101111101;
        12'd786: TDATA = 50'b01110011011001101110010000110111100101100101011100;
        12'd787: TDATA = 50'b01110011011000011010110100110111100011101100111000;
        12'd788: TDATA = 50'b01110011010111000111100100110111100001110100101001;
        12'd789: TDATA = 50'b01110011010101110100010000110111011111111100011001;
        12'd790: TDATA = 50'b01110011010100100001000000110111011110000100001111;
        12'd791: TDATA = 50'b01110011010011001101110110110111011100001100010000;
        12'd792: TDATA = 50'b01110011010001111010110000110111011010010100011001;
        12'd793: TDATA = 50'b01110011010000100111101000110111011000011100100100;
        12'd794: TDATA = 50'b01110011001111010100100010110111010110100100110011;
        12'd795: TDATA = 50'b01110011001110000001100100110111010100101101010000;
        12'd796: TDATA = 50'b01110011001100101110100110110111010010110101110001;
        12'd797: TDATA = 50'b01110011001011011011101010110111010000111110011000;
        12'd798: TDATA = 50'b01110011001010001000110010110111001111000111000110;
        12'd799: TDATA = 50'b01110011001000110101111110110111001101001111111100;
        12'd800: TDATA = 50'b01110011000111100011001100110111001011011000111000;
        12'd801: TDATA = 50'b01110011000110010000100000110111001001100010000000;
        12'd802: TDATA = 50'b01110011000100111101110000110111000111101011000110;
        12'd803: TDATA = 50'b01110011000011101011001000110111000101110100010111;
        12'd804: TDATA = 50'b01110011000010011000011100110111000011111101100111;
        12'd805: TDATA = 50'b01110011000001000101111000110111000010000111000110;
        12'd806: TDATA = 50'b01110010111111110011011000110111000000010000101101;
        12'd807: TDATA = 50'b01110010111110100000111000110110111110011010010110;
        12'd808: TDATA = 50'b01110010111101001110011100110110111100100100000101;
        12'd809: TDATA = 50'b01110010111011111100000010110110111010101101111100;
        12'd810: TDATA = 50'b01110010111010101001101110110110111000110111111110;
        12'd811: TDATA = 50'b01110010111001010111011010110110110111000010000011;
        12'd812: TDATA = 50'b01110010111000000101000110110110110101001100001010;
        12'd813: TDATA = 50'b01110010110110110010111010110110110011010110100001;
        12'd814: TDATA = 50'b01110010110101100000101010110110110001100000110010;
        12'd815: TDATA = 50'b01110010110100001110100010110110101111101011010011;
        12'd816: TDATA = 50'b01110010110010111100100000110110101101110101111110;
        12'd817: TDATA = 50'b01110010110001101010011010110110101100000000101000;
        12'd818: TDATA = 50'b01110010110000011000011100110110101010001011011101;
        12'd819: TDATA = 50'b01110010101111000110011010110110101000010110010001;
        12'd820: TDATA = 50'b01110010101101110100100000110110100110100001010100;
        12'd821: TDATA = 50'b01110010101100100010101010110110100100101100011110;
        12'd822: TDATA = 50'b01110010101011010000110010110110100010110111100110;
        12'd823: TDATA = 50'b01110010101001111111000010110110100001000010111101;
        12'd824: TDATA = 50'b01110010101000101101001110110110011111001110010011;
        12'd825: TDATA = 50'b01110010100111011011100010110110011101011001110100;
        12'd826: TDATA = 50'b01110010100110001001111000110110011011100101011100;
        12'd827: TDATA = 50'b01110010100100111000001110110110011001110001000111;
        12'd828: TDATA = 50'b01110010100011100110100110110110010111111100111000;
        12'd829: TDATA = 50'b01110010100010010101001000110110010110001000111001;
        12'd830: TDATA = 50'b01110010100001000011101010110110010100010100111100;
        12'd831: TDATA = 50'b01110010011111110010001010110110010010100000111110;
        12'd832: TDATA = 50'b01110010011110100000101110110110010000101101001011;
        12'd833: TDATA = 50'b01110010011101001111010110110110001110111001011110;
        12'd834: TDATA = 50'b01110010011011111110000010110110001101000101111001;
        12'd835: TDATA = 50'b01110010011010101100110000110110001011010010011010;
        12'd836: TDATA = 50'b01110010011001011011100000110110001001011111000010;
        12'd837: TDATA = 50'b01110010011000001010011000110110000111101011110101;
        12'd838: TDATA = 50'b01110010010110111001001100110110000101111000100111;
        12'd839: TDATA = 50'b01110010010101101000000010110110000100000101011111;
        12'd840: TDATA = 50'b01110010010100010111000000110110000010010010100011;
        12'd841: TDATA = 50'b01110010010011000101111010110110000000011111100100;
        12'd842: TDATA = 50'b01110010010001110101000000110101111110101100111010;
        12'd843: TDATA = 50'b01110010010000100100000000110101111100111010001001;
        12'd844: TDATA = 50'b01110010001111010011000110110101111011000111100011;
        12'd845: TDATA = 50'b01110010001110000010001110110101111001010101000100;
        12'd846: TDATA = 50'b01110010001100110001011010110101110111100010101100;
        12'd847: TDATA = 50'b01110010001011100000101010110101110101110000011011;
        12'd848: TDATA = 50'b01110010001010001111111000110101110011111110001100;
        12'd849: TDATA = 50'b01110010001000111111001110110101110010001100001000;
        12'd850: TDATA = 50'b01110010000111101110100010110101110000011010000111;
        12'd851: TDATA = 50'b01110010000110011101111110110101101110101000010000;
        12'd852: TDATA = 50'b01110010000101001101010110110101101100110110011000;
        12'd853: TDATA = 50'b01110010000011111100110100110101101011000100101011;
        12'd854: TDATA = 50'b01110010000010101100011000110101101001010011001001;
        12'd855: TDATA = 50'b01110010000001011011111000110101100111100001100101;
        12'd856: TDATA = 50'b01110010000000001011100010110101100101110000010001;
        12'd857: TDATA = 50'b01110001111110111011000110110101100011111110110110;
        12'd858: TDATA = 50'b01110001111101101010110100110101100010001101101011;
        12'd859: TDATA = 50'b01110001111100011010100000110101100000011100100010;
        12'd860: TDATA = 50'b01110001111011001010010000110101011110101011100000;
        12'd861: TDATA = 50'b01110001111001111010000100110101011100111010100100;
        12'd862: TDATA = 50'b01110001111000101001110110110101011011001001101011;
        12'd863: TDATA = 50'b01110001110111011001110110110101011001011001000101;
        12'd864: TDATA = 50'b01110001110110001001101110110101010111101000011010;
        12'd865: TDATA = 50'b01110001110100111001101110110101010101110111111001;
        12'd866: TDATA = 50'b01110001110011101001110000110101010100000111011111;
        12'd867: TDATA = 50'b01110001110010011001101110110101010010010111000011;
        12'd868: TDATA = 50'b01110001110001001001110100110101010000100110110010;
        12'd869: TDATA = 50'b01110001101111111001111100110101001110110110101000;
        12'd870: TDATA = 50'b01110001101110101010000110110101001101000110100101;
        12'd871: TDATA = 50'b01110001101101011010011000110101001011010110101100;
        12'd872: TDATA = 50'b01110001101100001010101000110101001001100110110110;
        12'd873: TDATA = 50'b01110001101010111010111010110101000111110111000010;
        12'd874: TDATA = 50'b01110001101001101011010000110101000110000111011001;
        12'd875: TDATA = 50'b01110001101000011011101010110101000100010111110111;
        12'd876: TDATA = 50'b01110001100111001100000010110101000010101000010011;
        12'd877: TDATA = 50'b01110001100101111100100010110101000000111000111110;
        12'd878: TDATA = 50'b01110001100100101100111110110100111111001001100111;
        12'd879: TDATA = 50'b01110001100011011101100010110100111101011010011100;
        12'd880: TDATA = 50'b01110001100010001110001000110100111011101011010110;
        12'd881: TDATA = 50'b01110001100000111110110000110100111001111100011000;
        12'd882: TDATA = 50'b01110001011111101111011010110100111000001101011100;
        12'd883: TDATA = 50'b01110001011110100000000110110100110110011110100110;
        12'd884: TDATA = 50'b01110001011101010000111000110100110100101111111011;
        12'd885: TDATA = 50'b01110001011100000001100110110100110011000001001111;
        12'd886: TDATA = 50'b01110001011010110010011110110100110001010010110001;
        12'd887: TDATA = 50'b01110001011001100011010110110100101111100100010110;
        12'd888: TDATA = 50'b01110001011000010100001110110100101101110101111101;
        12'd889: TDATA = 50'b01110001010111000101000110110100101100000111100111;
        12'd890: TDATA = 50'b01110001010101110110001010110100101010011001100100;
        12'd891: TDATA = 50'b01110001010100100111001100110100101000101011011111;
        12'd892: TDATA = 50'b01110001010011011000010010110100100110111101100100;
        12'd893: TDATA = 50'b01110001010010001001010110110100100101001111101000;
        12'd894: TDATA = 50'b01110001010000111010100000110100100011100001110111;
        12'd895: TDATA = 50'b01110001001111101011101110110100100001110100001100;
        12'd896: TDATA = 50'b01110001001110011100111110110100100000000110101000;
        12'd897: TDATA = 50'b01110001001101001110001110110100011110011001000110;
        12'd898: TDATA = 50'b01110001001011111111011110110100011100101011100111;
        12'd899: TDATA = 50'b01110001001010110000110110110100011010111110010110;
        12'd900: TDATA = 50'b01110001001001100010010000110100011001010001001000;
        12'd901: TDATA = 50'b01110001001000010011101100110100010111100100000001;
        12'd902: TDATA = 50'b01110001000111000101001010110100010101110110111111;
        12'd903: TDATA = 50'b01110001000101110110100110110100010100001001111101;
        12'd904: TDATA = 50'b01110001000100101000001100110100010010011101001001;
        12'd905: TDATA = 50'b01110001000011011001110100110100010000110000011011;
        12'd906: TDATA = 50'b01110001000010001011011100110100001111000011110000;
        12'd907: TDATA = 50'b01110001000000111101000100110100001101010111000111;
        12'd908: TDATA = 50'b01110000111111101110110010110100001011101010101001;
        12'd909: TDATA = 50'b01110000111110100000100000110100001001111110001101;
        12'd910: TDATA = 50'b01110000111101010010010100110100001000010001111100;
        12'd911: TDATA = 50'b01110000111100000100001000110100000110100101101101;
        12'd912: TDATA = 50'b01110000111010110101111110110100000100111001100101;
        12'd913: TDATA = 50'b01110000111001100111111000110100000011001101100011;
        12'd914: TDATA = 50'b01110000111000011001110110110100000001100001101000;
        12'd915: TDATA = 50'b01110000110111001011110110110011111111110101110011;
        12'd916: TDATA = 50'b01110000110101111101110110110011111110001010000000;
        12'd917: TDATA = 50'b01110000110100101111111000110011111100011110010100;
        12'd918: TDATA = 50'b01110000110011100001111110110011111010110010101111;
        12'd919: TDATA = 50'b01110000110010010100001010110011111001000111010100;
        12'd920: TDATA = 50'b01110000110001000110010110110011110111011011111011;
        12'd921: TDATA = 50'b01110000101111111000100110110011110101110000101001;
        12'd922: TDATA = 50'b01110000101110101010110010110011110100000101010101;
        12'd923: TDATA = 50'b01110000101101011101000110110011110010011010010000;
        12'd924: TDATA = 50'b01110000101100001111011110110011110000101111010001;
        12'd925: TDATA = 50'b01110000101011000001110110110011101111000100010100;
        12'd926: TDATA = 50'b01110000101001110100001110110011101101011001011010;
        12'd927: TDATA = 50'b01110000101000100110101010110011101011101110100110;
        12'd928: TDATA = 50'b01110000100111011001001110110011101010000100000001;
        12'd929: TDATA = 50'b01110000100110001011101110110011101000011001011010;
        12'd930: TDATA = 50'b01110000100100111110010010110011100110101110111001;
        12'd931: TDATA = 50'b01110000100011110000111010110011100101000100011111;
        12'd932: TDATA = 50'b01110000100010100011100100110011100011011010001011;
        12'd933: TDATA = 50'b01110000100001010110010000110011100001101111111110;
        12'd934: TDATA = 50'b01110000100000001001000000110011100000000101110111;
        12'd935: TDATA = 50'b01110000011110111011110000110011011110011011110010;
        12'd936: TDATA = 50'b01110000011101101110100000110011011100110001110000;
        12'd937: TDATA = 50'b01110000011100100001010110110011011011000111111000;
        12'd938: TDATA = 50'b01110000011011010100010010110011011001011110001011;
        12'd939: TDATA = 50'b01110000011010000111001110110011010111110100100000;
        12'd940: TDATA = 50'b01110000011000111010001010110011010110001010110111;
        12'd941: TDATA = 50'b01110000010111101101001010110011010100100001010100;
        12'd942: TDATA = 50'b01110000010110100000001100110011010010110111111000;
        12'd943: TDATA = 50'b01110000010101010011010100110011010001001110100110;
        12'd944: TDATA = 50'b01110000010100000110011100110011001111100101010111;
        12'd945: TDATA = 50'b01110000010010111001100100110011001101111100001010;
        12'd946: TDATA = 50'b01110000010001101100101110110011001100010011000011;
        12'd947: TDATA = 50'b01110000010000100000000000110011001010101010000111;
        12'd948: TDATA = 50'b01110000001111010011010000110011001001000001001100;
        12'd949: TDATA = 50'b01110000001110000110100010110011000111011000010101;
        12'd950: TDATA = 50'b01110000001100111001111000110011000101101111100111;
        12'd951: TDATA = 50'b01110000001011101101010010110011000100000111000000;
        12'd952: TDATA = 50'b01110000001010100000110000110011000010011110011111;
        12'd953: TDATA = 50'b01110000001001010100001010110011000000110101111101;
        12'd954: TDATA = 50'b01110000001000000111101010110010111111001101100101;
        12'd955: TDATA = 50'b01110000000110111011010000110010111101100101010111;
        12'd956: TDATA = 50'b01110000000101101110110010110010111011111101000111;
        12'd957: TDATA = 50'b01110000000100100010011000110010111010010100111110;
        12'd958: TDATA = 50'b01110000000011010110000010110010111000101100111011;
        12'd959: TDATA = 50'b01110000000010001001101110110010110111000100111110;
        12'd960: TDATA = 50'b01110000000000111101100000110010110101011101001011;
        12'd961: TDATA = 50'b01101111111111110001001110110010110011110101010111;
        12'd962: TDATA = 50'b01101111111110100101000000110010110010001101101001;
        12'd963: TDATA = 50'b01101111111101011000110110110010110000100110000010;
        12'd964: TDATA = 50'b01101111111100001100110000110010101110111110100100;
        12'd965: TDATA = 50'b01101111111011000000101100110010101101010111001001;
        12'd966: TDATA = 50'b01101111111001110100100110110010101011101111110000;
        12'd967: TDATA = 50'b01101111111000101000101010110010101010001000100110;
        12'd968: TDATA = 50'b01101111110111011100101100110010101000100001011001;
        12'd969: TDATA = 50'b01101111110110010000110010110010100110111010010111;
        12'd970: TDATA = 50'b01101111110101000100110100110010100101010011001111;
        12'd971: TDATA = 50'b01101111110011111001000000110010100011101100011010;
        12'd972: TDATA = 50'b01101111110010101101001010110010100010000101100010;
        12'd973: TDATA = 50'b01101111110001100001011000110010100000011110110001;
        12'd974: TDATA = 50'b01101111110000010101101000110010011110111000000110;
        12'd975: TDATA = 50'b01101111101111001001111110110010011101010001100101;
        12'd976: TDATA = 50'b01101111101101111110010000110010011011101011000011;
        12'd977: TDATA = 50'b01101111101100110010100110110010011010000100100111;
        12'd978: TDATA = 50'b01101111101011100111000110110010011000011110011001;
        12'd979: TDATA = 50'b01101111101010011011011110110010010110111000000101;
        12'd980: TDATA = 50'b01101111101001001111111110110010010101010001111011;
        12'd981: TDATA = 50'b01101111101000000100100010110010010011101011111100;
        12'd982: TDATA = 50'b01101111100110111001000010110010010010000101110110;
        12'd983: TDATA = 50'b01101111100101101101100110110010010000011111111011;
        12'd984: TDATA = 50'b01101111100100100010010010110010001110111010001010;
        12'd985: TDATA = 50'b01101111100011010111000000110010001101010100100000;
        12'd986: TDATA = 50'b01101111100010001011101010110010001011101110110011;
        12'd987: TDATA = 50'b01101111100001000000011000110010001010001001001101;
        12'd988: TDATA = 50'b01101111011111110101001010110010001000100011101101;
        12'd989: TDATA = 50'b01101111011110101010000000110010000110111110010111;
        12'd990: TDATA = 50'b01101111011101011110111000110010000101011001000011;
        12'd991: TDATA = 50'b01101111011100010011101110110010000011110011110010;
        12'd992: TDATA = 50'b01101111011011001000101100110010000010001110101010;
        12'd993: TDATA = 50'b01101111011001111101101000110010000000101001100101;
        12'd994: TDATA = 50'b01101111011000110010101000110001111111000100100110;
        12'd995: TDATA = 50'b01101111010111100111101100110001111101011111101101;
        12'd996: TDATA = 50'b01101111010110011100101110110001111011111010110110;
        12'd997: TDATA = 50'b01101111010101010001111000110001111010010110001001;
        12'd998: TDATA = 50'b01101111010100000111000000110001111000110001011111;
        12'd999: TDATA = 50'b01101111010010111100010000110001110111001100111111;
        12'd1000: TDATA = 50'b01101111010001110001011100110001110101101000011100;
        12'd1001: TDATA = 50'b01101111010000100110101110110001110100000100000100;
        12'd1002: TDATA = 50'b01101111001111011100000000110001110010011111101110;
        12'd1003: TDATA = 50'b01101111001110010001011000110001110000111011100010;
        12'd1004: TDATA = 50'b01101111001101000110110000110001101111010111011001;
        12'd1005: TDATA = 50'b01101111001011111100001000110001101101110011010001;
        12'd1006: TDATA = 50'b01101111001010110001100110110001101100001111010011;
        12'd1007: TDATA = 50'b01101111001001100111000100110001101010101011011000;
        12'd1008: TDATA = 50'b01101111001000011100100010110001101001000111011111;
        12'd1009: TDATA = 50'b01101111000111010010001000110001100111100011110100;
        12'd1010: TDATA = 50'b01101111000110000111110000110001100110000000001011;
        12'd1011: TDATA = 50'b01101111000100111101010100110001100100011100100000;
        12'd1012: TDATA = 50'b01101111000011110011000000110001100010111001000011;
        12'd1013: TDATA = 50'b01101111000010101000101110110001100001010101101000;
        12'd1014: TDATA = 50'b01101111000001011110011110110001011111110010010011;
        12'd1015: TDATA = 50'b01101111000000010100001110110001011110001111000001;
        12'd1016: TDATA = 50'b01101110111111001010000000110001011100101011110100;
        12'd1017: TDATA = 50'b01101110111101111111110110110001011011001000101110;
        12'd1018: TDATA = 50'b01101110111100110101110000110001011001100101101101;
        12'd1019: TDATA = 50'b01101110111011101011101100110001011000000010110011;
        12'd1020: TDATA = 50'b01101110111010100001101010110001010110011111111111;
        12'd1021: TDATA = 50'b01101110111001010111100110110001010100111101001001;
        12'd1022: TDATA = 50'b01101110111000001101101000110001010011011010011100;
        12'd1023: TDATA = 50'b01101110110111000011101010110001010001110111110010;
        12'd1024: TDATA = 50'b01101110110101111001110010110001010000010101010010;
        12'd1025: TDATA = 50'b01101110110100101111111010110001001110110010110101;
        12'd1026: TDATA = 50'b01101110110011100110000110110001001101010000011101;
        12'd1027: TDATA = 50'b01101110110010011100010100110001001011101110001011;
        12'd1028: TDATA = 50'b01101110110001010010100010110001001010001011111011;
        12'd1029: TDATA = 50'b01101110110000001000110110110001001000101001110101;
        12'd1030: TDATA = 50'b01101110101110111111001010110001000111000111110001;
        12'd1031: TDATA = 50'b01101110101101110101100000110001000101100101110100;
        12'd1032: TDATA = 50'b01101110101100101011111010110001000100000011111100;
        12'd1033: TDATA = 50'b01101110101011100010010010110001000010100010000010;
        12'd1034: TDATA = 50'b01101110101010011000110010110001000001000000010111;
        12'd1035: TDATA = 50'b01101110101001001111010010110000111111011110101101;
        12'd1036: TDATA = 50'b01101110101000000101110010110000111101111101000101;
        12'd1037: TDATA = 50'b01101110100110111100011000110000111100011011101000;
        12'd1038: TDATA = 50'b01101110100101110010111110110000111010111010001100;
        12'd1039: TDATA = 50'b01101110100100101001100110110000111001011000110111;
        12'd1040: TDATA = 50'b01101110100011100000010000110000110111110111100011;
        12'd1041: TDATA = 50'b01101110100010010110111110110000110110010110011001;
        12'd1042: TDATA = 50'b01101110100001001101101110110000110100110101010010;
        12'd1043: TDATA = 50'b01101110100000000100100000110000110011010100010000;
        12'd1044: TDATA = 50'b01101110011110111011010010110000110001110011010001;
        12'd1045: TDATA = 50'b01101110011101110010001010110000110000010010011011;
        12'd1046: TDATA = 50'b01101110011100101001000010110000101110110001101000;
        12'd1047: TDATA = 50'b01101110011011100000000000110000101101010000111110;
        12'd1048: TDATA = 50'b01101110011010010110111010110000101011110000010010;
        12'd1049: TDATA = 50'b01101110011001001101111100110000101010001111110000;
        12'd1050: TDATA = 50'b01101110011000000101000000110000101000101111010101;
        12'd1051: TDATA = 50'b01101110010110111100000000110000100111001110110111;
        12'd1052: TDATA = 50'b01101110010101110011001010110000100101101110100111;
        12'd1053: TDATA = 50'b01101110010100101010001110110000100100001110010001;
        12'd1054: TDATA = 50'b01101110010011100001011100110000100010101110001001;
        12'd1055: TDATA = 50'b01101110010010011000101000110000100001001110000011;
        12'd1056: TDATA = 50'b01101110010001001111110110110000011111101101111111;
        12'd1057: TDATA = 50'b01101110010000000111000110110000011110001110000001;
        12'd1058: TDATA = 50'b01101110001110111110011000110000011100101110001001;
        12'd1059: TDATA = 50'b01101110001101110101101110110000011011001110010111;
        12'd1060: TDATA = 50'b01101110001100101101001010110000011001101110101111;
        12'd1061: TDATA = 50'b01101110001011100100100100110000011000001111000101;
        12'd1062: TDATA = 50'b01101110001010011100000010110000010110101111100100;
        12'd1063: TDATA = 50'b01101110001001010011011110110000010101010000000010;
        12'd1064: TDATA = 50'b01101110001000001011000000110000010011110000101001;
        12'd1065: TDATA = 50'b01101110000111000010100110110000010010010001010111;
        12'd1066: TDATA = 50'b01101110000101111010001010110000010000110010000110;
        12'd1067: TDATA = 50'b01101110000100110001110010110000001111010010111011;
        12'd1068: TDATA = 50'b01101110000011101001011110110000001101110011110110;
        12'd1069: TDATA = 50'b01101110000010100001001100110000001100010100111000;
        12'd1070: TDATA = 50'b01101110000001011000110110110000001010110101110111;
        12'd1071: TDATA = 50'b01101110000000010000101000110000001001010111000000;
        12'd1072: TDATA = 50'b01101101111111001000011100110000000111111000001110;
        12'd1073: TDATA = 50'b01101101111110000000010010110000000110011001100011;
        12'd1074: TDATA = 50'b01101101111100111000001010110000000100111010111010;
        12'd1075: TDATA = 50'b01101101111011110000000000110000000011011100010010;
        12'd1076: TDATA = 50'b01101101111010101000000000110000000001111101111000;
        12'd1077: TDATA = 50'b01101101111001011111111110110000000000011111011101;
        12'd1078: TDATA = 50'b01101101111000010111111110101111111111000001000111;
        12'd1079: TDATA = 50'b01101101110111010000000000101111111101100010110111;
        12'd1080: TDATA = 50'b01101101110110001000000100101111111100000100101001;
        12'd1081: TDATA = 50'b01101101110101000000001010101111111010100110100000;
        12'd1082: TDATA = 50'b01101101110011111000010110101111111001001000100010;
        12'd1083: TDATA = 50'b01101101110010110000100010101111110111101010100101;
        12'd1084: TDATA = 50'b01101101110001101000101110101111110110001100101011;
        12'd1085: TDATA = 50'b01101101110000100000111010101111110100101110110010;
        12'd1086: TDATA = 50'b01101101101111011001001110101111110011010001000111;
        12'd1087: TDATA = 50'b01101101101110010001100100101111110001110011011110;
        12'd1088: TDATA = 50'b01101101101101001001111100101111110000010101111011;
        12'd1089: TDATA = 50'b01101101101100000010010100101111101110111000011001;
        12'd1090: TDATA = 50'b01101101101010111010101110101111101101011010111110;
        12'd1091: TDATA = 50'b01101101101001110011001010101111101011111101100100;
        12'd1092: TDATA = 50'b01101101101000101011101000101111101010100000010000;
        12'd1093: TDATA = 50'b01101101100111100100001100101111101001000011000110;
        12'd1094: TDATA = 50'b01101101100110011100110000101111100111100101111110;
        12'd1095: TDATA = 50'b01101101100101010101010100101111100110001000111000;
        12'd1096: TDATA = 50'b01101101100100001101111010101111100100101011110111;
        12'd1097: TDATA = 50'b01101101100011000110101000101111100011001111000001;
        12'd1098: TDATA = 50'b01101101100001111111010010101111100001110010001000;
        12'd1099: TDATA = 50'b01101101100000111000000010101111100000010101011001;
        12'd1100: TDATA = 50'b01101101011111110000110010101111011110111000101011;
        12'd1101: TDATA = 50'b01101101011110101001100010101111011101011100000000;
        12'd1102: TDATA = 50'b01101101011101100010011000101111011011111111011111;
        12'd1103: TDATA = 50'b01101101011100011011010000101111011010100011000011;
        12'd1104: TDATA = 50'b01101101011011010100001010101111011001000110101001;
        12'd1105: TDATA = 50'b01101101011010001101000110101111010111101010010100;
        12'd1106: TDATA = 50'b01101101011001000110000010101111010110001110000010;
        12'd1107: TDATA = 50'b01101101010111111111000100101111010100110001111001;
        12'd1108: TDATA = 50'b01101101010110111000000010101111010011010101101111;
        12'd1109: TDATA = 50'b01101101010101110001001000101111010001111001101110;
        12'd1110: TDATA = 50'b01101101010100101010010000101111010000011101110010;
        12'd1111: TDATA = 50'b01101101010011100011011000101111001111000001111001;
        12'd1112: TDATA = 50'b01101101010010011100100010101111001101100110000101;
        12'd1113: TDATA = 50'b01101101010001010101101110101111001100001010010011;
        12'd1114: TDATA = 50'b01101101010000001110111100101111001010101110100111;
        12'd1115: TDATA = 50'b01101101001111001000010000101111001001010011000101;
        12'd1116: TDATA = 50'b01101101001110000001100000101111000111110111100000;
        12'd1117: TDATA = 50'b01101101001100111010111000101111000110011100000101;
        12'd1118: TDATA = 50'b01101101001011110100001100101111000101000000101001;
        12'd1119: TDATA = 50'b01101101001010101101101000101111000011100101011001;
        12'd1120: TDATA = 50'b01101101001001100111000000101111000010001010000100;
        12'd1121: TDATA = 50'b01101101001000100000100000101111000000101110111100;
        12'd1122: TDATA = 50'b01101101000111011010000000101110111111010011110110;
        12'd1123: TDATA = 50'b01101101000110010011100110101110111101111000111010;
        12'd1124: TDATA = 50'b01101101000101001101000110101110111100011101110111;
        12'd1125: TDATA = 50'b01101101000100000110101110101110111011000011000010;
        12'd1126: TDATA = 50'b01101101000011000000010100101110111001101000001011;
        12'd1127: TDATA = 50'b01101101000001111001111110101110111000001101011010;
        12'd1128: TDATA = 50'b01101101000000110011101010101110110110110010101111;
        12'd1129: TDATA = 50'b01101100111111101101011100101110110101011000001101;
        12'd1130: TDATA = 50'b01101100111110100111001110101110110011111101101101;
        12'd1131: TDATA = 50'b01101100111101100001000000101110110010100011001110;
        12'd1132: TDATA = 50'b01101100111100011010111000101110110001001000111001;
        12'd1133: TDATA = 50'b01101100111011010100101010101110101111101110011111;
        12'd1134: TDATA = 50'b01101100111010001110101000101110101110010100010101;
        12'd1135: TDATA = 50'b01101100111001001000100010101110101100111010001010;
        12'd1136: TDATA = 50'b01101100111000000010011110101110101011100000000000;
        12'd1137: TDATA = 50'b01101100110110111100011110101110101010000110000000;
        12'd1138: TDATA = 50'b01101100110101110110100000101110101000101100000010;
        12'd1139: TDATA = 50'b01101100110100110000100110101110100111010010001101;
        12'd1140: TDATA = 50'b01101100110011101010101010101110100101111000010110;
        12'd1141: TDATA = 50'b01101100110010100100110010101110100100011110100101;
        12'd1142: TDATA = 50'b01101100110001011110111110101110100011000100111101;
        12'd1143: TDATA = 50'b01101100110000011001001100101110100001101011010111;
        12'd1144: TDATA = 50'b01101100101111010011010110101110100000010001101111;
        12'd1145: TDATA = 50'b01101100101110001101101100101110011110111000011001;
        12'd1146: TDATA = 50'b01101100101101000111111100101110011101011110111100;
        12'd1147: TDATA = 50'b01101100101100000010001110101110011100000101100101;
        12'd1148: TDATA = 50'b01101100101010111100101000101110011010101100011000;
        12'd1149: TDATA = 50'b01101100101001110111000100101110011001010011010000;
        12'd1150: TDATA = 50'b01101100101000110001011100101110010111111010000110;
        12'd1151: TDATA = 50'b01101100100111101011111000101110010110100001000001;
        12'd1152: TDATA = 50'b01101100100110100110011000101110010101001000000011;
        12'd1153: TDATA = 50'b01101100100101100000111010101110010011101111001001;
        12'd1154: TDATA = 50'b01101100100100011011011110101110010010010110010110;
        12'd1155: TDATA = 50'b01101100100011010110000100101110010000111101100100;
        12'd1156: TDATA = 50'b01101100100010010000101100101110001111100100111000;
        12'd1157: TDATA = 50'b01101100100001001011010100101110001110001100001110;
        12'd1158: TDATA = 50'b01101100100000000101111110101110001100110011101001;
        12'd1159: TDATA = 50'b01101100011111000000110000101110001011011011001110;
        12'd1160: TDATA = 50'b01101100011101111011011110101110001010000010110000;
        12'd1161: TDATA = 50'b01101100011100110110001110101110001000101010011001;
        12'd1162: TDATA = 50'b01101100011011110001000010101110000111010010000110;
        12'd1163: TDATA = 50'b01101100011010101011111010101110000101111001111010;
        12'd1164: TDATA = 50'b01101100011001100110110100101110000100100001110011;
        12'd1165: TDATA = 50'b01101100011000100001101110101110000011001001101110;
        12'd1166: TDATA = 50'b01101100010111011100101000101110000001110001101010;
        12'd1167: TDATA = 50'b01101100010110010111101000101110000000011001110000;
        12'd1168: TDATA = 50'b01101100010101010010101000101101111111000001111000;
        12'd1169: TDATA = 50'b01101100010100001101101000101101111101101010000001;
        12'd1170: TDATA = 50'b01101100010011001000101110101101111100010010010100;
        12'd1171: TDATA = 50'b01101100010010000011110100101101111010111010101000;
        12'd1172: TDATA = 50'b01101100010000111110111100101101111001100011000010;
        12'd1173: TDATA = 50'b01101100001111111010000110101101111000001011011110;
        12'd1174: TDATA = 50'b01101100001110110101010010101101110110110100000000;
        12'd1175: TDATA = 50'b01101100001101110000100100101101110101011100101010;
        12'd1176: TDATA = 50'b01101100001100101011110110101101110100000101010111;
        12'd1177: TDATA = 50'b01101100001011100111001000101101110010101110000101;
        12'd1178: TDATA = 50'b01101100001010100010011010101101110001010110110101;
        12'd1179: TDATA = 50'b01101100001001011101110010101101101111111111101110;
        12'd1180: TDATA = 50'b01101100001000011001001100101101101110101000101101;
        12'd1181: TDATA = 50'b01101100000111010100101000101101101101010001101110;
        12'd1182: TDATA = 50'b01101100000110010000000110101101101011111010110100;
        12'd1183: TDATA = 50'b01101100000101001011100100101101101010100011111011;
        12'd1184: TDATA = 50'b01101100000100000111000100101101101001001101001001;
        12'd1185: TDATA = 50'b01101100000011000010100110101101100111110110011000;
        12'd1186: TDATA = 50'b01101100000001111110001100101101100110011111110000;
        12'd1187: TDATA = 50'b01101100000000111001110110101101100101001001001110;
        12'd1188: TDATA = 50'b01101011111111110101011110101101100011110010101010;
        12'd1189: TDATA = 50'b01101011111110110001001010101101100010011100001111;
        12'd1190: TDATA = 50'b01101011111101101100111000101101100001000101110110;
        12'd1191: TDATA = 50'b01101011111100101000101000101101011111101111100010;
        12'd1192: TDATA = 50'b01101011111011100100011000101101011110011001010000;
        12'd1193: TDATA = 50'b01101011111010100000001010101101011101000011000011;
        12'd1194: TDATA = 50'b01101011111001011100000000101101011011101100111100;
        12'd1195: TDATA = 50'b01101011111000010111110110101101011010010110110111;
        12'd1196: TDATA = 50'b01101011110111010011110000101101011001000000110111;
        12'd1197: TDATA = 50'b01101011110110001111101100101101010111101010111101;
        12'd1198: TDATA = 50'b01101011110101001011101010101101010110010101001000;
        12'd1199: TDATA = 50'b01101011110100000111101010101101010100111111010101;
        12'd1200: TDATA = 50'b01101011110011000011101100101101010011101001100111;
        12'd1201: TDATA = 50'b01101011110001111111101110101101010010010011111011;
        12'd1202: TDATA = 50'b01101011110000111011110010101101010000111110010100;
        12'd1203: TDATA = 50'b01101011101111110111111010101101001111101000110011;
        12'd1204: TDATA = 50'b01101011101110110100000010101101001110010011010100;
        12'd1205: TDATA = 50'b01101011101101110000010000101101001100111101111110;
        12'd1206: TDATA = 50'b01101011101100101100011110101101001011101000101001;
        12'd1207: TDATA = 50'b01101011101011101000110000101101001010010011011010;
        12'd1208: TDATA = 50'b01101011101010100100111110101101001000111110001001;
        12'd1209: TDATA = 50'b01101011101001100001010010101101000111101001000001;
        12'd1210: TDATA = 50'b01101011101000011101101000101101000110010011111111;
        12'd1211: TDATA = 50'b01101011100111011010000000101101000100111110111110;
        12'd1212: TDATA = 50'b01101011100110010110011100101101000011101010000110;
        12'd1213: TDATA = 50'b01101011100101010010110100101101000010010101001001;
        12'd1214: TDATA = 50'b01101011100100001111010100101101000001000000011000;
        12'd1215: TDATA = 50'b01101011100011001011110000101100111111101011100110;
        12'd1216: TDATA = 50'b01101011100010001000010100101100111110010110111100;
        12'd1217: TDATA = 50'b01101011100001000100111010101100111101000010011000;
        12'd1218: TDATA = 50'b01101011100000000001011010101100111011101101101110;
        12'd1219: TDATA = 50'b01101011011110111110000110101100111010011001010101;
        12'd1220: TDATA = 50'b01101011011101111010101110101100111001000100111010;
        12'd1221: TDATA = 50'b01101011011100110111011000101100110111110000100000;
        12'd1222: TDATA = 50'b01101011011011110100000110101100110110011100010000;
        12'd1223: TDATA = 50'b01101011011010110000110110101100110101001000000001;
        12'd1224: TDATA = 50'b01101011011001101101101000101100110011110011111000;
        12'd1225: TDATA = 50'b01101011011000101010011010101100110010011111110000;
        12'd1226: TDATA = 50'b01101011010111100111001110101100110001001011101110;
        12'd1227: TDATA = 50'b01101011010110100100000110101100101111110111110001;
        12'd1228: TDATA = 50'b01101011010101100000111110101100101110100011110101;
        12'd1229: TDATA = 50'b01101011010100011101111010101100101101001111111111;
        12'd1230: TDATA = 50'b01101011010011011010111000101100101011111100001111;
        12'd1231: TDATA = 50'b01101011010010010111110110101100101010101000100000;
        12'd1232: TDATA = 50'b01101011010001010100110110101100101001010100110110;
        12'd1233: TDATA = 50'b01101011010000010001111010101100101000000001010010;
        12'd1234: TDATA = 50'b01101011001111001110111110101100100110101101110000;
        12'd1235: TDATA = 50'b01101011001110001100000110101100100101011010010011;
        12'd1236: TDATA = 50'b01101011001101001001010010101100100100000110111111;
        12'd1237: TDATA = 50'b01101011001100000110011010101100100010110011100101;
        12'd1238: TDATA = 50'b01101011001011000011100110101100100001100000010100;
        12'd1239: TDATA = 50'b01101011001010000000110110101100100000001101001001;
        12'd1240: TDATA = 50'b01101011001000111110000110101100011110111001111111;
        12'd1241: TDATA = 50'b01101011000111111011010110101100011101100110110110;
        12'd1242: TDATA = 50'b01101011000110111000110000101100011100010011111011;
        12'd1243: TDATA = 50'b01101011000101110110000010101100011011000000111010;
        12'd1244: TDATA = 50'b01101011000100110011011100101100011001101110000010;
        12'd1245: TDATA = 50'b01101011000011110000111000101100011000011011001111;
        12'd1246: TDATA = 50'b01101011000010101110010100101100010111001000011110;
        12'd1247: TDATA = 50'b01101011000001101011110000101100010101110101101110;
        12'd1248: TDATA = 50'b01101011000000101001010010101100010100100011001000;
        12'd1249: TDATA = 50'b01101010111111100110110100101100010011010000100011;
        12'd1250: TDATA = 50'b01101010111110100100010110101100010001111101111111;
        12'd1251: TDATA = 50'b01101010111101100001111110101100010000101011100101;
        12'd1252: TDATA = 50'b01101010111100011111100110101100001111011001001100;
        12'd1253: TDATA = 50'b01101010111011011101001110101100001110000110110101;
        12'd1254: TDATA = 50'b01101010111010011010111100101100001100110100100111;
        12'd1255: TDATA = 50'b01101010111001011000101010101100001011100010011011;
        12'd1256: TDATA = 50'b01101010111000010110011000101100001010010000010000;
        12'd1257: TDATA = 50'b01101010110111010100001100101100001000111110001110;
        12'd1258: TDATA = 50'b01101010110110010010000000101100000111101100001110;
        12'd1259: TDATA = 50'b01101010110101001111110100101100000110011010001111;
        12'd1260: TDATA = 50'b01101010110100001101101010101100000101001000010110;
        12'd1261: TDATA = 50'b01101010110011001011100100101100000011110110100010;
        12'd1262: TDATA = 50'b01101010110010001001011110101100000010100100110000;
        12'd1263: TDATA = 50'b01101010110001000111011100101100000001010011000010;
        12'd1264: TDATA = 50'b01101010110000000101011100101100000000000001011010;
        12'd1265: TDATA = 50'b01101010101111000011011100101011111110101111110100;
        12'd1266: TDATA = 50'b01101010101110000001100010101011111101011110010111;
        12'd1267: TDATA = 50'b01101010101100111111100010101011111100001100110100;
        12'd1268: TDATA = 50'b01101010101011111101101010101011111010111011011101;
        12'd1269: TDATA = 50'b01101010101010111011110100101011111001101010001000;
        12'd1270: TDATA = 50'b01101010101001111001111100101011111000011000110101;
        12'd1271: TDATA = 50'b01101010101000111000001100101011110111000111101011;
        12'd1272: TDATA = 50'b01101010100111110110011000101011110101110110011110;
        12'd1273: TDATA = 50'b01101010100110110100101010101011110100100101011011;
        12'd1274: TDATA = 50'b01101010100101110010111100101011110011010100011001;
        12'd1275: TDATA = 50'b01101010100100110001001110101011110010000011011000;
        12'd1276: TDATA = 50'b01101010100011101111100010101011110000110010011101;
        12'd1277: TDATA = 50'b01101010100010101101111010101011101111100001100111;
        12'd1278: TDATA = 50'b01101010100001101100010110101011101110010000110111;
        12'd1279: TDATA = 50'b01101010100000101010110000101011101101000000000111;
        12'd1280: TDATA = 50'b01101010011111101001001110101011101011101111011110;
        12'd1281: TDATA = 50'b01101010011110100111110000101011101010011110111001;
        12'd1282: TDATA = 50'b01101010011101100110001110101011101001001110010010;
        12'd1283: TDATA = 50'b01101010011100100100110010101011100111111101110101;
        12'd1284: TDATA = 50'b01101010011011100011010110101011100110101101011000;
        12'd1285: TDATA = 50'b01101010011010100010000000101011100101011101000101;
        12'd1286: TDATA = 50'b01101010011001100000100110101011100100001100101111;
        12'd1287: TDATA = 50'b01101010011000011111010100101011100010111100100011;
        12'd1288: TDATA = 50'b01101010010111011101111110101011100001101100010100;
        12'd1289: TDATA = 50'b01101010010110011100101110101011100000011100001110;
        12'd1290: TDATA = 50'b01101010010101011011011110101011011111001100001010;
        12'd1291: TDATA = 50'b01101010010100011010001110101011011101111100000111;
        12'd1292: TDATA = 50'b01101010010011011001000100101011011100101100001101;
        12'd1293: TDATA = 50'b01101010010010010111110110101011011011011100010001;
        12'd1294: TDATA = 50'b01101010010001010110110000101011011010001100011110;
        12'd1295: TDATA = 50'b01101010010000010101101100101011011000111100110000;
        12'd1296: TDATA = 50'b01101010001111010100101000101011010111101101000100;
        12'd1297: TDATA = 50'b01101010001110010011100100101011010110011101011001;
        12'd1298: TDATA = 50'b01101010001101010010100010101011010101001101110011;
        12'd1299: TDATA = 50'b01101010001100010001100010101011010011111110001111;
        12'd1300: TDATA = 50'b01101010001011010000100110101011010010101110110100;
        12'd1301: TDATA = 50'b01101010001010001111101100101011010001011111011010;
        12'd1302: TDATA = 50'b01101010001001001110110100101011010000010000000101;
        12'd1303: TDATA = 50'b01101010001000001101111100101011001111000000110010;
        12'd1304: TDATA = 50'b01101010000111001101000110101011001101110001100100;
        12'd1305: TDATA = 50'b01101010000110001100010010101011001100100010011000;
        12'd1306: TDATA = 50'b01101010000101001011100000101011001011010011010001;
        12'd1307: TDATA = 50'b01101010000100001010101110101011001010000100001011;
        12'd1308: TDATA = 50'b01101010000011001010000010101011001000110101001110;
        12'd1309: TDATA = 50'b01101010000010001001010110101011000111100110010011;
        12'd1310: TDATA = 50'b01101010000001001000101100101011000110010111011101;
        12'd1311: TDATA = 50'b01101010000000001000000100101011000101001000101000;
        12'd1312: TDATA = 50'b01101001111111000111011010101011000011111001110101;
        12'd1313: TDATA = 50'b01101001111110000110111000101011000010101011001010;
        12'd1314: TDATA = 50'b01101001111101000110010100101011000001011100100001;
        12'd1315: TDATA = 50'b01101001111100000101110010101011000000001101111010;
        12'd1316: TDATA = 50'b01101001111011000101010010101010111110111111011000;
        12'd1317: TDATA = 50'b01101001111010000100110100101010111101110000111011;
        12'd1318: TDATA = 50'b01101001111001000100011000101010111100100010011111;
        12'd1319: TDATA = 50'b01101001111000000011111110101010111011010100001001;
        12'd1320: TDATA = 50'b01101001110111000011101010101010111010000101111011;
        12'd1321: TDATA = 50'b01101001110110000011010000101010111000110111101000;
        12'd1322: TDATA = 50'b01101001110101000010111100101010110111101001011101;
        12'd1323: TDATA = 50'b01101001110100000010101010101010110110011011010111;
        12'd1324: TDATA = 50'b01101001110011000010011010101010110101001101010011;
        12'd1325: TDATA = 50'b01101001110010000010001100101010110011111111010100;
        12'd1326: TDATA = 50'b01101001110001000001111110101010110010110001010111;
        12'd1327: TDATA = 50'b01101001110000000001110010101010110001100011011110;
        12'd1328: TDATA = 50'b01101001101111000001101010101010110000010101101011;
        12'd1329: TDATA = 50'b01101001101110000001100010101010101111000111111001;
        12'd1330: TDATA = 50'b01101001101101000001011010101010101101111010001001;
        12'd1331: TDATA = 50'b01101001101100000001010110101010101100101100011110;
        12'd1332: TDATA = 50'b01101001101011000001010100101010101011011110111000;
        12'd1333: TDATA = 50'b01101001101010000001010100101010101010010001010111;
        12'd1334: TDATA = 50'b01101001101001000001010110101010101001000011110111;
        12'd1335: TDATA = 50'b01101001101000000001011010101010100111110110011101;
        12'd1336: TDATA = 50'b01101001100111000001011110101010100110101001000100;
        12'd1337: TDATA = 50'b01101001100110000001100100101010100101011011110000;
        12'd1338: TDATA = 50'b01101001100101000001101110101010100100001110100001;
        12'd1339: TDATA = 50'b01101001100100000001111000101010100011000001010100;
        12'd1340: TDATA = 50'b01101001100011000010000110101010100001110100001100;
        12'd1341: TDATA = 50'b01101001100010000010010010101010100000100111000101;
        12'd1342: TDATA = 50'b01101001100001000010100010101010011111011010000011;
        12'd1343: TDATA = 50'b01101001100000000010110110101010011110001101000110;
        12'd1344: TDATA = 50'b01101001011111000011001100101010011101000000001111;
        12'd1345: TDATA = 50'b01101001011110000011011110101010011011110011010101;
        12'd1346: TDATA = 50'b01101001011101000011111000101010011010100110100100;
        12'd1347: TDATA = 50'b01101001011100000100001110101010011001011001110001;
        12'd1348: TDATA = 50'b01101001011011000100101010101010011000001101000110;
        12'd1349: TDATA = 50'b01101001011010000101000110101010010111000000011101;
        12'd1350: TDATA = 50'b01101001011001000101100100101010010101110011111001;
        12'd1351: TDATA = 50'b01101001011000000110000100101010010100100111010111;
        12'd1352: TDATA = 50'b01101001010111000110100110101010010011011010111001;
        12'd1353: TDATA = 50'b01101001010110000111001010101010010010001110100001;
        12'd1354: TDATA = 50'b01101001010101000111110000101010010001000010001010;
        12'd1355: TDATA = 50'b01101001010100001000011000101010001111110101111000;
        12'd1356: TDATA = 50'b01101001010011001001000010101010001110101001101011;
        12'd1357: TDATA = 50'b01101001010010001001101010101010001101011101011100;
        12'd1358: TDATA = 50'b01101001010001001010011000101010001100010001010101;
        12'd1359: TDATA = 50'b01101001010000001011000110101010001011000101010000;
        12'd1360: TDATA = 50'b01101001001111001011111000101010001001111001010000;
        12'd1361: TDATA = 50'b01101001001110001100101100101010001000101101010101;
        12'd1362: TDATA = 50'b01101001001101001101011100101010000111100001011000;
        12'd1363: TDATA = 50'b01101001001100001110010100101010000110010101100100;
        12'd1364: TDATA = 50'b01101001001011001111001000101010000101001001101101;
        12'd1365: TDATA = 50'b01101001001010010000000100101010000011111110000010;
        12'd1366: TDATA = 50'b01101001001001010000111100101010000010110010010010;
        12'd1367: TDATA = 50'b01101001001000010001111100101010000001100110101110;
        12'd1368: TDATA = 50'b01101001000111010010111000101010000000011011001000;
        12'd1369: TDATA = 50'b01101001000110010011111000101001111111001111100111;
        12'd1370: TDATA = 50'b01101001000101010100111000101001111110000100000111;
        12'd1371: TDATA = 50'b01101001000100010110000010101001111100111000110011;
        12'd1372: TDATA = 50'b01101001000011010111000010101001111011101101010110;
        12'd1373: TDATA = 50'b01101001000010011000001110101001111010100010001001;
        12'd1374: TDATA = 50'b01101001000001011001010100101001111001010110110110;
        12'd1375: TDATA = 50'b01101001000000011010100000101001111000001011101100;
        12'd1376: TDATA = 50'b01101000111111011011101100101001110111000000100011;
        12'd1377: TDATA = 50'b01101000111110011100111010101001110101110101011111;
        12'd1378: TDATA = 50'b01101000111101011110001010101001110100101010011100;
        12'd1379: TDATA = 50'b01101000111100011111011110101001110011011111100010;
        12'd1380: TDATA = 50'b01101000111011100000101110101001110010010100100010;
        12'd1381: TDATA = 50'b01101000111010100010000110101001110001001001101111;
        12'd1382: TDATA = 50'b01101000111001100011011010101001101111111110111001;
        12'd1383: TDATA = 50'b01101000111000100100110110101001101110110100001100;
        12'd1384: TDATA = 50'b01101000110111100110010000101001101101101001100000;
        12'd1385: TDATA = 50'b01101000110110100111101100101001101100011110110101;
        12'd1386: TDATA = 50'b01101000110101101001001010101001101011010100010000;
        12'd1387: TDATA = 50'b01101000110100101010101010101001101010001001101111;
        12'd1388: TDATA = 50'b01101000110011101100001100101001101000111111010000;
        12'd1389: TDATA = 50'b01101000110010101101110000101001100111110100110110;
        12'd1390: TDATA = 50'b01101000110001101111010110101001100110101010100001;
        12'd1391: TDATA = 50'b01101000110000110000111010101001100101100000001001;
        12'd1392: TDATA = 50'b01101000101111110010100010101001100100010101110111;
        12'd1393: TDATA = 50'b01101000101110110100001110101001100011001011101101;
        12'd1394: TDATA = 50'b01101000101101110101111100101001100010000001100100;
        12'd1395: TDATA = 50'b01101000101100110111100110101001100000110111011010;
        12'd1396: TDATA = 50'b01101000101011111001010110101001011111101101011000;
        12'd1397: TDATA = 50'b01101000101010111011001100101001011110100011011110;
        12'd1398: TDATA = 50'b01101000101001111100111100101001011101011001011110;
        12'd1399: TDATA = 50'b01101000101000111110101110101001011100001111100100;
        12'd1400: TDATA = 50'b01101000101000000000101000101001011011000101110010;
        12'd1401: TDATA = 50'b01101000100111000010100000101001011001111100000001;
        12'd1402: TDATA = 50'b01101000100110000100011010101001011000110010010010;
        12'd1403: TDATA = 50'b01101000100101000110010110101001010111101000100111;
        12'd1404: TDATA = 50'b01101000100100001000010010101001010110011110111110;
        12'd1405: TDATA = 50'b01101000100011001010010100101001010101010101011110;
        12'd1406: TDATA = 50'b01101000100010001100010010101001010100001011111011;
        12'd1407: TDATA = 50'b01101000100001001110010100101001010011000010011101;
        12'd1408: TDATA = 50'b01101000100000010000011010101001010001111001000100;
        12'd1409: TDATA = 50'b01101000011111010010011110101001010000101111101101;
        12'd1410: TDATA = 50'b01101000011110010100100110101001001111100110011010;
        12'd1411: TDATA = 50'b01101000011101010110101110101001001110011101001001;
        12'd1412: TDATA = 50'b01101000011100011000111100101001001101010100000000;
        12'd1413: TDATA = 50'b01101000011011011011001010101001001100001010111001;
        12'd1414: TDATA = 50'b01101000011010011101011000101001001011000001110011;
        12'd1415: TDATA = 50'b01101000011001011111100110101001001001111000101110;
        12'd1416: TDATA = 50'b01101000011000100001111000101001001000101111101110;
        12'd1417: TDATA = 50'b01101000010111100100001100101001000111100110110011;
        12'd1418: TDATA = 50'b01101000010110100110100010101001000110011101111101;
        12'd1419: TDATA = 50'b01101000010101101000111100101001000101010101001100;
        12'd1420: TDATA = 50'b01101000010100101011010100101001000100001100011001;
        12'd1421: TDATA = 50'b01101000010011101101110000101001000011000011101110;
        12'd1422: TDATA = 50'b01101000010010110000001000101001000001111010111101;
        12'd1423: TDATA = 50'b01101000010001110010101000101001000000110010011000;
        12'd1424: TDATA = 50'b01101000010000110101001000101000111111101001110101;
        12'd1425: TDATA = 50'b01101000001111110111101000101000111110100001010011;
        12'd1426: TDATA = 50'b01101000001110111010001110101000111101011000111001;
        12'd1427: TDATA = 50'b01101000001101111100110000101000111100010000011101;
        12'd1428: TDATA = 50'b01101000001100111111011010101000111011001000001010;
        12'd1429: TDATA = 50'b01101000001100000010000000101000111001111111110100;
        12'd1430: TDATA = 50'b01101000001011000100101000101000111000110111100011;
        12'd1431: TDATA = 50'b01101000001010000111010100101000110111101111010111;
        12'd1432: TDATA = 50'b01101000001001001010000100101000110110100111010000;
        12'd1433: TDATA = 50'b01101000001000001100110010101000110101011111001011;
        12'd1434: TDATA = 50'b01101000000111001111100010101000110100010111000110;
        12'd1435: TDATA = 50'b01101000000110010010010100101000110011001111000111;
        12'd1436: TDATA = 50'b01101000000101010101000110101000110010000111001000;
        12'd1437: TDATA = 50'b01101000000100010111111110101000110000111111010010;
        12'd1438: TDATA = 50'b01101000000011011010110010101000101111110111011010;
        12'd1439: TDATA = 50'b01101000000010011101101110101000101110101111101011;
        12'd1440: TDATA = 50'b01101000000001100000101000101000101101100111111100;
        12'd1441: TDATA = 50'b01101000000000100011100110101000101100100000010011;
        12'd1442: TDATA = 50'b01100111111111100110100100101000101011011000101011;
        12'd1443: TDATA = 50'b01100111111110101001100010101000101010010001000100;
        12'd1444: TDATA = 50'b01100111111101101100100100101000101001001001100010;
        12'd1445: TDATA = 50'b01100111111100101111101000101000101000000010000100;
        12'd1446: TDATA = 50'b01100111111011110010101110101000100110111010101100;
        12'd1447: TDATA = 50'b01100111111010110101110010101000100101110011010001;
        12'd1448: TDATA = 50'b01100111111001111000111010101000100100101011111011;
        12'd1449: TDATA = 50'b01100111111000111100000110101000100011100100101110;
        12'd1450: TDATA = 50'b01100111110111111111001110101000100010011101011011;
        12'd1451: TDATA = 50'b01100111110111000010011110101000100001010110010011;
        12'd1452: TDATA = 50'b01100111110110000101101110101000100000001111001101;
        12'd1453: TDATA = 50'b01100111110101001000111110101000011111001000001001;
        12'd1454: TDATA = 50'b01100111110100001100001110101000011110000001000101;
        12'd1455: TDATA = 50'b01100111110011001111100100101000011100111010001010;
        12'd1456: TDATA = 50'b01100111110010010010110110101000011011110011001101;
        12'd1457: TDATA = 50'b01100111110001010110010000101000011010101100010111;
        12'd1458: TDATA = 50'b01100111110000011001101000101000011001100101100100;
        12'd1459: TDATA = 50'b01100111101111011101000010101000011000011110110001;
        12'd1460: TDATA = 50'b01100111101110100000011110101000010111011000000011;
        12'd1461: TDATA = 50'b01100111101101100011111100101000010110010001011011;
        12'd1462: TDATA = 50'b01100111101100100111011100101000010101001010110011;
        12'd1463: TDATA = 50'b01100111101011101010111110101000010100000100010000;
        12'd1464: TDATA = 50'b01100111101010101110100000101000010010111101101111;
        12'd1465: TDATA = 50'b01100111101001110010000010101000010001110111001110;
        12'd1466: TDATA = 50'b01100111101000110101101010101000010000110000110110;
        12'd1467: TDATA = 50'b01100111100111111001010010101000001111101010100000;
        12'd1468: TDATA = 50'b01100111100110111100111010101000001110100100001010;
        12'd1469: TDATA = 50'b01100111100110000000101000101000001101011101111101;
        12'd1470: TDATA = 50'b01100111100101000100010010101000001100010111101110;
        12'd1471: TDATA = 50'b01100111100100001000000100101000001011010001100111;
        12'd1472: TDATA = 50'b01100111100011001011110010101000001010001011011101;
        12'd1473: TDATA = 50'b01100111100010001111100010101000001001000101011001;
        12'd1474: TDATA = 50'b01100111100001010011010100101000000111111111010110;
        12'd1475: TDATA = 50'b01100111100000010111001000101000000110111001010111;
        12'd1476: TDATA = 50'b01100111011111011011000010101000000101110011100001;
        12'd1477: TDATA = 50'b01100111011110011110111100101000000100101101101100;
        12'd1478: TDATA = 50'b01100111011101100010110010101000000011100111110101;
        12'd1479: TDATA = 50'b01100111011100100110110000101000000010100010000110;
        12'd1480: TDATA = 50'b01100111011011101010101100101000000001011100011000;
        12'd1481: TDATA = 50'b01100111011010101110101010101000000000010110101100;
        12'd1482: TDATA = 50'b01100111011001110010101010100111111111010001000100;
        12'd1483: TDATA = 50'b01100111011000110110101100100111111110001011100001;
        12'd1484: TDATA = 50'b01100111010111111010101100100111111101000101111100;
        12'd1485: TDATA = 50'b01100111010110111110110110100111111100000000100010;
        12'd1486: TDATA = 50'b01100111010110000010111000100111111010111011000011;
        12'd1487: TDATA = 50'b01100111010101000111000010100111111001110101101100;
        12'd1488: TDATA = 50'b01100111010100001011001110100111111000110000011010;
        12'd1489: TDATA = 50'b01100111010011001111011010100111110111101011001001;
        12'd1490: TDATA = 50'b01100111010010010011100110100111110110100101111001;
        12'd1491: TDATA = 50'b01100111010001010111111000100111110101100000110001;
        12'd1492: TDATA = 50'b01100111010000011100000110100111110100011011101000;
        12'd1493: TDATA = 50'b01100111001111100000011000100111110011010110100011;
        12'd1494: TDATA = 50'b01100111001110100100101010100111110010010001011111;
        12'd1495: TDATA = 50'b01100111001101101001000010100111110001001100100011;
        12'd1496: TDATA = 50'b01100111001100101101011010100111110000000111101001;
        12'd1497: TDATA = 50'b01100111001011110001110010100111101111000010110000;
        12'd1498: TDATA = 50'b01100111001010110110001010100111101101111101111000;
        12'd1499: TDATA = 50'b01100111001001111010101000100111101100111001001000;
        12'd1500: TDATA = 50'b01100111001000111111000100100111101011110100010110;
        12'd1501: TDATA = 50'b01100111001000000011100100100111101010101111101101;
        12'd1502: TDATA = 50'b01100111000111001000000110100111101001101011000100;
        12'd1503: TDATA = 50'b01100111000110001100100110100111101000100110011101;
        12'd1504: TDATA = 50'b01100111000101010001001010100111100111100001111010;
        12'd1505: TDATA = 50'b01100111000100010101110010100111100110011101011100;
        12'd1506: TDATA = 50'b01100111000011011010010110100111100101011000111100;
        12'd1507: TDATA = 50'b01100111000010011111000010100111100100010100101000;
        12'd1508: TDATA = 50'b01100111000001100011101010100111100011010000001101;
        12'd1509: TDATA = 50'b01100111000000101000010110100111100010001011111011;
        12'd1510: TDATA = 50'b01100110111111101101000100100111100001000111101010;
        12'd1511: TDATA = 50'b01100110111110110001110100100111100000000011011110;
        12'd1512: TDATA = 50'b01100110111101110110100100100111011110111111010011;
        12'd1513: TDATA = 50'b01100110111100111011010110100111011101111011001101;
        12'd1514: TDATA = 50'b01100110111100000000001010100111011100110111001000;
        12'd1515: TDATA = 50'b01100110111011000101000000100111011011110011001000;
        12'd1516: TDATA = 50'b01100110111010001001110110100111011010101111001001;
        12'd1517: TDATA = 50'b01100110111001001110101110100111011001101011001110;
        12'd1518: TDATA = 50'b01100110111000010011101010100111011000100111011000;
        12'd1519: TDATA = 50'b01100110110111011000100110100111010111100011100100;
        12'd1520: TDATA = 50'b01100110110110011101100010100111010110011111110000;
        12'd1521: TDATA = 50'b01100110110101100010100010100111010101011100000010;
        12'd1522: TDATA = 50'b01100110110100100111100100100111010100011000011000;
        12'd1523: TDATA = 50'b01100110110011101100100110100111010011010100101111;
        12'd1524: TDATA = 50'b01100110110010110001101010100111010010010001001011;
        12'd1525: TDATA = 50'b01100110110001110110110000100111010001001101101000;
        12'd1526: TDATA = 50'b01100110110000111011111000100111010000001010001001;
        12'd1527: TDATA = 50'b01100110110000000001000000100111001111000110101100;
        12'd1528: TDATA = 50'b01100110101111000110001000100111001110000011010000;
        12'd1529: TDATA = 50'b01100110101110001011010010100111001100111111111001;
        12'd1530: TDATA = 50'b01100110101101010000100000100111001011111100100110;
        12'd1531: TDATA = 50'b01100110101100010101101110100111001010111001010101;
        12'd1532: TDATA = 50'b01100110101011011011000000100111001001110110001000;
        12'd1533: TDATA = 50'b01100110101010100000010100100111001000110011000000;
        12'd1534: TDATA = 50'b01100110101001100101101000100111000111101111111001;
        12'd1535: TDATA = 50'b01100110101000101010111100100111000110101100110011;
        12'd1536: TDATA = 50'b01100110100111110000010000100111000101101001101111;
        12'd1537: TDATA = 50'b01100110100110110101101100100111000100100110110101;
        12'd1538: TDATA = 50'b01100110100101111011000100100111000011100011110111;
        12'd1539: TDATA = 50'b01100110100101000000100000100111000010100001000000;
        12'd1540: TDATA = 50'b01100110100100000101111110100111000001011110001010;
        12'd1541: TDATA = 50'b01100110100011001011011110100111000000011011011010;
        12'd1542: TDATA = 50'b01100110100010010000111110100110111111011000101010;
        12'd1543: TDATA = 50'b01100110100001010110011110100110111110010101111011;
        12'd1544: TDATA = 50'b01100110100000011011111110100110111101010011001110;
        12'd1545: TDATA = 50'b01100110011111100001100100100110111100010000101001;
        12'd1546: TDATA = 50'b01100110011110100111001010100110111011001110000101;
        12'd1547: TDATA = 50'b01100110011101101100110110100110111010001011101001;
        12'd1548: TDATA = 50'b01100110011100110010011100100110111001001001000111;
        12'd1549: TDATA = 50'b01100110011011111000001000100110111000000110101101;
        12'd1550: TDATA = 50'b01100110011010111101110100100110110111000100010100;
        12'd1551: TDATA = 50'b01100110011010000011100010100110110110000010000001;
        12'd1552: TDATA = 50'b01100110011001001001010010100110110100111111101110;
        12'd1553: TDATA = 50'b01100110011000001111000100100110110011111101100000;
        12'd1554: TDATA = 50'b01100110010111010100110110100110110010111011010011;
        12'd1555: TDATA = 50'b01100110010110011010101010100110110001111001001010;
        12'd1556: TDATA = 50'b01100110010101100000100010100110110000110111000110;
        12'd1557: TDATA = 50'b01100110010100100110011010100110101111110101000100;
        12'd1558: TDATA = 50'b01100110010011101100010010100110101110110011000010;
        12'd1559: TDATA = 50'b01100110010010110010001010100110101101110001000010;
        12'd1560: TDATA = 50'b01100110010001111000001000100110101100101111001010;
        12'd1561: TDATA = 50'b01100110010000111110000110100110101011101101010010;
        12'd1562: TDATA = 50'b01100110010000000100000100100110101010101011011100;
        12'd1563: TDATA = 50'b01100110001111001010000110100110101001101001101011;
        12'd1564: TDATA = 50'b01100110001110010000000110100110101000100111111011;
        12'd1565: TDATA = 50'b01100110001101010110001010100110100111100110001111;
        12'd1566: TDATA = 50'b01100110001100011100010010100110100110100100101000;
        12'd1567: TDATA = 50'b01100110001011100010010110100110100101100010111110;
        12'd1568: TDATA = 50'b01100110001010101000100010100110100100100001100001;
        12'd1569: TDATA = 50'b01100110001001101110101010100110100011011111111101;
        12'd1570: TDATA = 50'b01100110001000110100110110100110100010011110100001;
        12'd1571: TDATA = 50'b01100110000111111011000100100110100001011101000111;
        12'd1572: TDATA = 50'b01100110000111000001010100100110100000011011110001;
        12'd1573: TDATA = 50'b01100110000110000111100100100110011111011010011100;
        12'd1574: TDATA = 50'b01100110000101001101110100100110011110011001001000;
        12'd1575: TDATA = 50'b01100110000100010100000110100110011101010111111001;
        12'd1576: TDATA = 50'b01100110000011011010011010100110011100010110101011;
        12'd1577: TDATA = 50'b01100110000010100000110010100110011011010101100101;
        12'd1578: TDATA = 50'b01100110000001100111001100100110011010010100100000;
        12'd1579: TDATA = 50'b01100110000000101101100010100110011001010011011001;
        12'd1580: TDATA = 50'b01100101111111110011111110100110011000010010011010;
        12'd1581: TDATA = 50'b01100101111110111010011010100110010111010001011100;
        12'd1582: TDATA = 50'b01100101111110000000111000100110010110010000100010;
        12'd1583: TDATA = 50'b01100101111101000111011000100110010101001111101010;
        12'd1584: TDATA = 50'b01100101111100001101110110100110010100001110110010;
        12'd1585: TDATA = 50'b01100101111011010100011100100110010011001110000011;
        12'd1586: TDATA = 50'b01100101111010011010111110100110010010001101010001;
        12'd1587: TDATA = 50'b01100101111001100001100010100110010001001100100100;
        12'd1588: TDATA = 50'b01100101111000101000001010100110010000001011111100;
        12'd1589: TDATA = 50'b01100101110111101110110010100110001111001011010100;
        12'd1590: TDATA = 50'b01100101110110110101011010100110001110001010101110;
        12'd1591: TDATA = 50'b01100101110101111100001000100110001101001010010000;
        12'd1592: TDATA = 50'b01100101110101000010110110100110001100001001110010;
        12'd1593: TDATA = 50'b01100101110100001001100100100110001011001001010110;
        12'd1594: TDATA = 50'b01100101110011010000010010100110001010001000111011;
        12'd1595: TDATA = 50'b01100101110010010111000100100110001001001000100101;
        12'd1596: TDATA = 50'b01100101110001011101111000100110001000001000010011;
        12'd1597: TDATA = 50'b01100101110000100100101100100110000111001000000010;
        12'd1598: TDATA = 50'b01100101101111101011100010100110000110000111110110;
        12'd1599: TDATA = 50'b01100101101110110010011100100110000101000111101110;
        12'd1600: TDATA = 50'b01100101101101111001010100100110000100000111100100;
        12'd1601: TDATA = 50'b01100101101101000000010000100110000011000111100001;
        12'd1602: TDATA = 50'b01100101101100000111001000100110000010000111011010;
        12'd1603: TDATA = 50'b01100101101011001110001000100110000001000111011101;
        12'd1604: TDATA = 50'b01100101101010010101001000100110000000000111100001;
        12'd1605: TDATA = 50'b01100101101001011100001000100101111111000111100111;
        12'd1606: TDATA = 50'b01100101101000100011001000100101111110000111101110;
        12'd1607: TDATA = 50'b01100101100111101010001110100101111101000111111100;
        12'd1608: TDATA = 50'b01100101100110110001010000100101111100001000001001;
        12'd1609: TDATA = 50'b01100101100101111000011010100101111011001000011101;
        12'd1610: TDATA = 50'b01100101100100111111100010100101111010001000110010;
        12'd1611: TDATA = 50'b01100101100100000110101000100101111001001001000101;
        12'd1612: TDATA = 50'b01100101100011001101110100100101111000001001100000;
        12'd1613: TDATA = 50'b01100101100010010101000100100101110111001001111111;
        12'd1614: TDATA = 50'b01100101100001011100010000100101110110001010011100;
        12'd1615: TDATA = 50'b01100101100000100011100010100101110101001011000001;
        12'd1616: TDATA = 50'b01100101011111101010110000100101110100001011100100;
        12'd1617: TDATA = 50'b01100101011110110010000010100101110011001100001011;
        12'd1618: TDATA = 50'b01100101011101111001011000100101110010001100110111;
        12'd1619: TDATA = 50'b01100101011101000000101100100101110001001101100011;
        12'd1620: TDATA = 50'b01100101011100001000000010100101110000001110010001;
        12'd1621: TDATA = 50'b01100101011011001111011010100101101111001111000011;
        12'd1622: TDATA = 50'b01100101011010010110111000100101101110001111111101;
        12'd1623: TDATA = 50'b01100101011001011110010010100101101101010000110101;
        12'd1624: TDATA = 50'b01100101011000100101101110100101101100010001101110;
        12'd1625: TDATA = 50'b01100101010111101101001100100101101011010010101011;
        12'd1626: TDATA = 50'b01100101010110110100101100100101101010010011101101;
        12'd1627: TDATA = 50'b01100101010101111100001110100101101001010100110000;
        12'd1628: TDATA = 50'b01100101010101000011110010100101101000010101110111;
        12'd1629: TDATA = 50'b01100101010100001011010110100101100111010111000000;
        12'd1630: TDATA = 50'b01100101010011010010111010100101100110011000001001;
        12'd1631: TDATA = 50'b01100101010010011010100000100101100101011001010111;
        12'd1632: TDATA = 50'b01100101010001100010001010100101100100011010101001;
        12'd1633: TDATA = 50'b01100101010000101001110010100101100011011011111010;
        12'd1634: TDATA = 50'b01100101001111110001100010100101100010011101010101;
        12'd1635: TDATA = 50'b01100101001110111001001110100101100001011110101110;
        12'd1636: TDATA = 50'b01100101001110000000111100100101100000100000001000;
        12'd1637: TDATA = 50'b01100101001101001000101100100101011111100001100110;
        12'd1638: TDATA = 50'b01100101001100010000011100100101011110100011000110;
        12'd1639: TDATA = 50'b01100101001011011000001110100101011101100100101010;
        12'd1640: TDATA = 50'b01100101001010100000000010100101011100100110001111;
        12'd1641: TDATA = 50'b01100101001001100111111010100101011011100111111100;
        12'd1642: TDATA = 50'b01100101001000101111110100100101011010101001101010;
        12'd1643: TDATA = 50'b01100101000111110111101010100101011001101011010101;
        12'd1644: TDATA = 50'b01100101000110111111100010100101011000101101000101;
        12'd1645: TDATA = 50'b01100101000110000111011110100101010111101110111010;
        12'd1646: TDATA = 50'b01100101000101001111011110100101010110110000110011;
        12'd1647: TDATA = 50'b01100101000100010111011010100101010101110010101001;
        12'd1648: TDATA = 50'b01100101000011011111011100100101010100110100101000;
        12'd1649: TDATA = 50'b01100101000010100111011110100101010011110110100111;
        12'd1650: TDATA = 50'b01100101000001101111100000100101010010111000100111;
        12'd1651: TDATA = 50'b01100101000000110111100010100101010001111010101001;
        12'd1652: TDATA = 50'b01100100111111111111101010100101010000111100110010;
        12'd1653: TDATA = 50'b01100100111111000111101110100101001111111110111001;
        12'd1654: TDATA = 50'b01100100111110001111111010100101001111000001001000;
        12'd1655: TDATA = 50'b01100100111101011000000100100101001110000011011000;
        12'd1656: TDATA = 50'b01100100111100100000010000100101001101000101101001;
        12'd1657: TDATA = 50'b01100100111011101000011110100101001100000111111110;
        12'd1658: TDATA = 50'b01100100111010110000101100100101001011001010010100;
        12'd1659: TDATA = 50'b01100100111001111000111010100101001010001100101100;
        12'd1660: TDATA = 50'b01100100111001000001001110100101001001001111001011;
        12'd1661: TDATA = 50'b01100100111000001001011110100101001000010001101000;
        12'd1662: TDATA = 50'b01100100110111010001110010100101000111010100001001;
        12'd1663: TDATA = 50'b01100100110110011010001010100101000110010110101110;
        12'd1664: TDATA = 50'b01100100110101100010100100100101000101011001011000;
        12'd1665: TDATA = 50'b01100100110100101010111000100101000100011011111101;
        12'd1666: TDATA = 50'b01100100110011110011010100100101000011011110101100;
        12'd1667: TDATA = 50'b01100100110010111011101110100101000010100001011001;
        12'd1668: TDATA = 50'b01100100110010000100001100100101000001100100001010;
        12'd1669: TDATA = 50'b01100100110001001100101100100101000000100111000000;
        12'd1670: TDATA = 50'b01100100110000010101001100100100111111101001110111;
        12'd1671: TDATA = 50'b01100100101111011101101100100100111110101100101111;
        12'd1672: TDATA = 50'b01100100101110100110001110100100111101101111101011;
        12'd1673: TDATA = 50'b01100100101101101110110010100100111100110010101001;
        12'd1674: TDATA = 50'b01100100101100110111010100100100111011110101100111;
        12'd1675: TDATA = 50'b01100100101011111111111110100100111010111000101101;
        12'd1676: TDATA = 50'b01100100101011001000101010100100111001111011111000;
        12'd1677: TDATA = 50'b01100100101010010001010010100100111000111111000000;
        12'd1678: TDATA = 50'b01100100101001011001111100100100111000000010001001;
        12'd1679: TDATA = 50'b01100100101000100010101000100100110111000101010110;
        12'd1680: TDATA = 50'b01100100100111101011010110100100110110001000101000;
        12'd1681: TDATA = 50'b01100100100110110100000110100100110101001011111011;
        12'd1682: TDATA = 50'b01100100100101111100111000100100110100001111010010;
        12'd1683: TDATA = 50'b01100100100101000101101010100100110011010010101011;
        12'd1684: TDATA = 50'b01100100100100001110011110100100110010010110000111;
        12'd1685: TDATA = 50'b01100100100011010111010100100100110001011001100101;
        12'd1686: TDATA = 50'b01100100100010100000001100100100110000011101000111;
        12'd1687: TDATA = 50'b01100100100001101001000100100100101111100000101010;
        12'd1688: TDATA = 50'b01100100100000110001111100100100101110100100001110;
        12'd1689: TDATA = 50'b01100100011111111010110110100100101101100111110110;
        12'd1690: TDATA = 50'b01100100011111000011110010100100101100101011100000;
        12'd1691: TDATA = 50'b01100100011110001100110000100100101011101111001101;
        12'd1692: TDATA = 50'b01100100011101010101101110100100101010110010111100;
        12'd1693: TDATA = 50'b01100100011100011110101110100100101001110110101111;
        12'd1694: TDATA = 50'b01100100011011100111110000100100101000111010100011;
        12'd1695: TDATA = 50'b01100100011010110000110100100100100111111110011100;
        12'd1696: TDATA = 50'b01100100011001111001111010100100100111000010011000;
        12'd1697: TDATA = 50'b01100100011001000010111110100100100110000110010011;
        12'd1698: TDATA = 50'b01100100011000001100000110100100100101001010010010;
        12'd1699: TDATA = 50'b01100100010111010101010010100100100100001110011000;
        12'd1700: TDATA = 50'b01100100010110011110011010100100100011010010011001;
        12'd1701: TDATA = 50'b01100100010101100111100110100100100010010110100001;
        12'd1702: TDATA = 50'b01100100010100110000110100100100100001011010101011;
        12'd1703: TDATA = 50'b01100100010011111010000100100100100000011110111000;
        12'd1704: TDATA = 50'b01100100010011000011010100100100011111100011000111;
        12'd1705: TDATA = 50'b01100100010010001100100100100100011110100111010111;
        12'd1706: TDATA = 50'b01100100010001010101110110100100011101101011101011;
        12'd1707: TDATA = 50'b01100100010000011111001010100100011100110000000000;
        12'd1708: TDATA = 50'b01100100001111101000100000100100011011110100011001;
        12'd1709: TDATA = 50'b01100100001110110001110110100100011010111000110100;
        12'd1710: TDATA = 50'b01100100001101111011001110100100011001111101010010;
        12'd1711: TDATA = 50'b01100100001101000100101000100100011001000001110010;
        12'd1712: TDATA = 50'b01100100001100001110000100100100011000000110010110;
        12'd1713: TDATA = 50'b01100100001011010111100000100100010111001010111011;
        12'd1714: TDATA = 50'b01100100001010100000111110100100010110001111100100;
        12'd1715: TDATA = 50'b01100100001001101010011110100100010101010100001110;
        12'd1716: TDATA = 50'b01100100001000110100000000100100010100011000111101;
        12'd1717: TDATA = 50'b01100100000111111101100010100100010011011101101100;
        12'd1718: TDATA = 50'b01100100000111000111000100100100010010100010011101;
        12'd1719: TDATA = 50'b01100100000110010000101000100100010001100111010010;
        12'd1720: TDATA = 50'b01100100000101011010001110100100010000101100001000;
        12'd1721: TDATA = 50'b01100100000100100011110110100100001111110001000010;
        12'd1722: TDATA = 50'b01100100000011101101011110100100001110110101111101;
        12'd1723: TDATA = 50'b01100100000010110111001100100100001101111010111111;
        12'd1724: TDATA = 50'b01100100000010000000110110100100001101000000000000;
        12'd1725: TDATA = 50'b01100100000001001010100100100100001100000101000100;
        12'd1726: TDATA = 50'b01100100000000010100010010100100001011001010001010;
        12'd1727: TDATA = 50'b01100011111111011110000100100100001010001111010100;
        12'd1728: TDATA = 50'b01100011111110100111110010100100001001010100011011;
        12'd1729: TDATA = 50'b01100011111101110001100110100100001000011001101010;
        12'd1730: TDATA = 50'b01100011111100111011011010100100000111011110111010;
        12'd1731: TDATA = 50'b01100011111100000101010000100100000110100100001111;
        12'd1732: TDATA = 50'b01100011111011001111001000100100000101101001100100;
        12'd1733: TDATA = 50'b01100011111010011000111100100100000100101110110111;
        12'd1734: TDATA = 50'b01100011111001100010111000100100000011110100010101;
        12'd1735: TDATA = 50'b01100011111000101100110010100100000010111001110001;
        12'd1736: TDATA = 50'b01100011110111110110110000100100000001111111010000;
        12'd1737: TDATA = 50'b01100011110111000000101100100100000001000100110001;
        12'd1738: TDATA = 50'b01100011110110001010101100100100000000001010010110;
        12'd1739: TDATA = 50'b01100011110101010100101100100011111111001111111100;
        12'd1740: TDATA = 50'b01100011110100011110101100100011111110010101100011;
        12'd1741: TDATA = 50'b01100011110011101000110010100011111101011011010010;
        12'd1742: TDATA = 50'b01100011110010110010110110100011111100100000111110;
        12'd1743: TDATA = 50'b01100011110001111100111100100011111011100110101110;
        12'd1744: TDATA = 50'b01100011110001000111000010100011111010101100100000;
        12'd1745: TDATA = 50'b01100011110000010001001110100011111001110010011001;
        12'd1746: TDATA = 50'b01100011101111011011010110100011111000111000001111;
        12'd1747: TDATA = 50'b01100011101110100101100010100011110111111110001010;
        12'd1748: TDATA = 50'b01100011101101101111101110100011110111000100000110;
        12'd1749: TDATA = 50'b01100011101100111001111110100011110110001010000110;
        12'd1750: TDATA = 50'b01100011101100000100001010100011110101010000000100;
        12'd1751: TDATA = 50'b01100011101011001110011100100011110100010110001001;
        12'd1752: TDATA = 50'b01100011101010011000101110100011110011011100001111;
        12'd1753: TDATA = 50'b01100011101001100011000010100011110010100010011010;
        12'd1754: TDATA = 50'b01100011101000101101011000100011110001101000100101;
        12'd1755: TDATA = 50'b01100011100111110111110000100011110000101110110101;
        12'd1756: TDATA = 50'b01100011100111000010001000100011101111110101000101;
        12'd1757: TDATA = 50'b01100011100110001100100000100011101110111011010111;
        12'd1758: TDATA = 50'b01100011100101010110111000100011101110000001101001;
        12'd1759: TDATA = 50'b01100011100100100001010010100011101101001000000000;
        12'd1760: TDATA = 50'b01100011100011101011110000100011101100001110011011;
        12'd1761: TDATA = 50'b01100011100010110110001110100011101011010100110111;
        12'd1762: TDATA = 50'b01100011100010000000110000100011101010011011010111;
        12'd1763: TDATA = 50'b01100011100001001011001110100011101001100001110100;
        12'd1764: TDATA = 50'b01100011100000010101110010100011101000101000011010;
        12'd1765: TDATA = 50'b01100011011111100000010110100011100111101111000000;
        12'd1766: TDATA = 50'b01100011011110101010111010100011100110110101100111;
        12'd1767: TDATA = 50'b01100011011101110101100000100011100101111100010010;
        12'd1768: TDATA = 50'b01100011011101000000001010100011100101000011000010;
        12'd1769: TDATA = 50'b01100011011100001010110010100011100100001001101111;
        12'd1770: TDATA = 50'b01100011011011010101011110100011100011010000100100;
        12'd1771: TDATA = 50'b01100011011010100000000110100011100010010111010011;
        12'd1772: TDATA = 50'b01100011011001101010110110100011100001011110001100;
        12'd1773: TDATA = 50'b01100011011000110101100110100011100000100101000111;
        12'd1774: TDATA = 50'b01100011011000000000010010100011011111101100000000;
        12'd1775: TDATA = 50'b01100011010111001011000110100011011110110011000000;
        12'd1776: TDATA = 50'b01100011010110010101110110100011011101111001111101;
        12'd1777: TDATA = 50'b01100011010101100000101100100011011101000001000010;
        12'd1778: TDATA = 50'b01100011010100101011011110100011011100001000000101;
        12'd1779: TDATA = 50'b01100011010011110110011000100011011011001111001111;
        12'd1780: TDATA = 50'b01100011010011000001001110100011011010010110010111;
        12'd1781: TDATA = 50'b01100011010010001100000110100011011001011101100011;
        12'd1782: TDATA = 50'b01100011010001010111000010100011011000100100110011;
        12'd1783: TDATA = 50'b01100011010000100001111110100011010111101100000100;
        12'd1784: TDATA = 50'b01100011001111101100111010100011010110110011010110;
        12'd1785: TDATA = 50'b01100011001110110111111010100011010101111010101100;
        12'd1786: TDATA = 50'b01100011001110000010111000100011010101000010000011;
        12'd1787: TDATA = 50'b01100011001101001101111010100011010100001001011111;
        12'd1788: TDATA = 50'b01100011001100011000111100100011010011010000111011;
        12'd1789: TDATA = 50'b01100011001011100011111110100011010010011000011000;
        12'd1790: TDATA = 50'b01100011001010101111000110100011010001011111111100;
        12'd1791: TDATA = 50'b01100011001001111010001110100011010000100111100010;
        12'd1792: TDATA = 50'b01100011001001000101010110100011001111101111001000;
        12'd1793: TDATA = 50'b01100011001000010000011110100011001110110110110000;
        12'd1794: TDATA = 50'b01100011000111011011100110100011001101111110011000;
        12'd1795: TDATA = 50'b01100011000110100110110010100011001101000110000100;
        12'd1796: TDATA = 50'b01100011000101110010000000100011001100001101110101;
        12'd1797: TDATA = 50'b01100011000100111101001110100011001011010101100111;
        12'd1798: TDATA = 50'b01100011000100001000011110100011001010011101011100;
        12'd1799: TDATA = 50'b01100011000011010011110000100011001001100101010011;
        12'd1800: TDATA = 50'b01100011000010011111000100100011001000101101001101;
        12'd1801: TDATA = 50'b01100011000001101010011000100011000111110101001001;
        12'd1802: TDATA = 50'b01100011000000110101101100100011000110111101000101;
        12'd1803: TDATA = 50'b01100011000000000001000000100011000110000101000011;
        12'd1804: TDATA = 50'b01100010111111001100010110100011000101001101000101;
        12'd1805: TDATA = 50'b01100010111110010111110000100011000100010101001010;
        12'd1806: TDATA = 50'b01100010111101100011001000100011000011011101001110;
        12'd1807: TDATA = 50'b01100010111100101110101000100011000010100101011100;
        12'd1808: TDATA = 50'b01100010111011111010000100100011000001101101100111;
        12'd1809: TDATA = 50'b01100010111011000101100010100011000000110101110100;
        12'd1810: TDATA = 50'b01100010111010010001000010100010111111111110000101;
        12'd1811: TDATA = 50'b01100010111001011100100010100010111111000110010110;
        12'd1812: TDATA = 50'b01100010111000101000000010100010111110001110101001;
        12'd1813: TDATA = 50'b01100010110111110011100100100010111101010111000000;
        12'd1814: TDATA = 50'b01100010110110111111001110100010111100011111011101;
        12'd1815: TDATA = 50'b01100010110110001010110000100010111011100111110110;
        12'd1816: TDATA = 50'b01100010110101010110011010100010111010110000010110;
        12'd1817: TDATA = 50'b01100010110100100010000000100010111001111000110011;
        12'd1818: TDATA = 50'b01100010110011101101101000100010111001000001010101;
        12'd1819: TDATA = 50'b01100010110010111001010100100010111000001001111011;
        12'd1820: TDATA = 50'b01100010110010000101000100100010110111010010100101;
        12'd1821: TDATA = 50'b01100010110001010000110000100010110110011011001100;
        12'd1822: TDATA = 50'b01100010110000011100011110100010110101100011111000;
        12'd1823: TDATA = 50'b01100010101111101000001110100010110100101100100100;
        12'd1824: TDATA = 50'b01100010101110110100000010100010110011110101011000;
        12'd1825: TDATA = 50'b01100010101101111111110010100010110010111110000111;
        12'd1826: TDATA = 50'b01100010101101001011100110100010110010000110111100;
        12'd1827: TDATA = 50'b01100010101100010111011110100010110001001111110110;
        12'd1828: TDATA = 50'b01100010101011100011010110100010110000011000110001;
        12'd1829: TDATA = 50'b01100010101010101111001110100010101111100001101100;
        12'd1830: TDATA = 50'b01100010101001111011000110100010101110101010101001;
        12'd1831: TDATA = 50'b01100010101001000110111110100010101101110011100110;
        12'd1832: TDATA = 50'b01100010101000010010111100100010101100111100101011;
        12'd1833: TDATA = 50'b01100010100111011110111010100010101100000101110000;
        12'd1834: TDATA = 50'b01100010100110101010111000100010101011001110110111;
        12'd1835: TDATA = 50'b01100010100101110110110110100010101010010111111110;
        12'd1836: TDATA = 50'b01100010100101000010111000100010101001100001001001;
        12'd1837: TDATA = 50'b01100010100100001110111100100010101000101010011001;
        12'd1838: TDATA = 50'b01100010100011011011000000100010100111110011101001;
        12'd1839: TDATA = 50'b01100010100010100111000100100010100110111100111011;
        12'd1840: TDATA = 50'b01100010100001110011001010100010100110000110010000;
        12'd1841: TDATA = 50'b01100010100000111111010010100010100101001111100110;
        12'd1842: TDATA = 50'b01100010100000001011011100100010100100011001000000;
        12'd1843: TDATA = 50'b01100010011111010111100110100010100011100010011100;
        12'd1844: TDATA = 50'b01100010011110100011110000100010100010101011111000;
        12'd1845: TDATA = 50'b01100010011101101111111010100010100001110101010101;
        12'd1846: TDATA = 50'b01100010011100111100001010100010100000111110111001;
        12'd1847: TDATA = 50'b01100010011100001000011010100010100000001000011110;
        12'd1848: TDATA = 50'b01100010011011010100101010100010011111010010000100;
        12'd1849: TDATA = 50'b01100010011010100000111010100010011110011011101011;
        12'd1850: TDATA = 50'b01100010011001101101010000100010011101100101011001;
        12'd1851: TDATA = 50'b01100010011000111001100010100010011100101111000101;
        12'd1852: TDATA = 50'b01100010011000000101111000100010011011111000110100;
        12'd1853: TDATA = 50'b01100010010111010010001110100010011011000010100101;
        12'd1854: TDATA = 50'b01100010010110011110101000100010011010001100011010;
        12'd1855: TDATA = 50'b01100010010101101011000000100010011001010110010000;
        12'd1856: TDATA = 50'b01100010010100110111011010100010011000100000000110;
        12'd1857: TDATA = 50'b01100010010100000011110110100010010111101010000001;
        12'd1858: TDATA = 50'b01100010010011010000010100100010010110110011111111;
        12'd1859: TDATA = 50'b01100010010010011100110100100010010101111101111111;
        12'd1860: TDATA = 50'b01100010010001101001010010100010010101000111111111;
        12'd1861: TDATA = 50'b01100010010000110101110010100010010100010010000001;
        12'd1862: TDATA = 50'b01100010010000000010010100100010010011011100000110;
        12'd1863: TDATA = 50'b01100010001111001110111000100010010010100110001111;
        12'd1864: TDATA = 50'b01100010001110011011011110100010010001110000011010;
        12'd1865: TDATA = 50'b01100010001101101000000010100010010000111010100101;
        12'd1866: TDATA = 50'b01100010001100110100101010100010010000000100110100;
        12'd1867: TDATA = 50'b01100010001100000001010010100010001111001111000100;
        12'd1868: TDATA = 50'b01100010001011001101111010100010001110011001010100;
        12'd1869: TDATA = 50'b01100010001010011010101000100010001101100011101101;
        12'd1870: TDATA = 50'b01100010001001100111010100100010001100101110000010;
        12'd1871: TDATA = 50'b01100010001000110100000010100010001011111000011100;
        12'd1872: TDATA = 50'b01100010001000000000110000100010001011000010110111;
        12'd1873: TDATA = 50'b01100010000111001101100100100010001010001101011000;
        12'd1874: TDATA = 50'b01100010000110011010010010100010001001010111110101;
        12'd1875: TDATA = 50'b01100010000101100111000110100010001000100010011000;
        12'd1876: TDATA = 50'b01100010000100110011111010100010000111101100111101;
        12'd1877: TDATA = 50'b01100010000100000000101110100010000110110111100010;
        12'd1878: TDATA = 50'b01100010000011001101100100100010000110000010001011;
        12'd1879: TDATA = 50'b01100010000010011010011100100010000101001100110101;
        12'd1880: TDATA = 50'b01100010000001100111010010100010000100010111100001;
        12'd1881: TDATA = 50'b01100010000000110100010000100010000011100010010011;
        12'd1882: TDATA = 50'b01100010000000000001001010100010000010101101000011;
        12'd1883: TDATA = 50'b01100001111111001110000100100010000001110111110011;
        12'd1884: TDATA = 50'b01100001111110011011000100100010000001000010101011;
        12'd1885: TDATA = 50'b01100001111101101000000100100010000000001101100100;
        12'd1886: TDATA = 50'b01100001111100110101000100100001111111011000011101;
        12'd1887: TDATA = 50'b01100001111100000010000100100001111110100011011000;
        12'd1888: TDATA = 50'b01100001111011001111001010100001111101101110011001;
        12'd1889: TDATA = 50'b01100001111010011100001010100001111100111001010110;
        12'd1890: TDATA = 50'b01100001111001101001010000100001111100000100011001;
        12'd1891: TDATA = 50'b01100001111000110110010110100001111011001111011101;
        12'd1892: TDATA = 50'b01100001111000000011100010100001111010011010101000;
        12'd1893: TDATA = 50'b01100001110111010000101000100001111001100101101110;
        12'd1894: TDATA = 50'b01100001110110011101110000100001111000110000111000;
        12'd1895: TDATA = 50'b01100001110101101010111100100001110111111100000110;
        12'd1896: TDATA = 50'b01100001110100111000001100100001110111000111011000;
        12'd1897: TDATA = 50'b01100001110100000101011000100001110110010010100111;
        12'd1898: TDATA = 50'b01100001110011010010101010100001110101011101111110;
        12'd1899: TDATA = 50'b01100001110010011111110110100001110100101001001111;
        12'd1900: TDATA = 50'b01100001110001101101001010100001110011110100101010;
        12'd1901: TDATA = 50'b01100001110000111010011100100001110011000000000100;
        12'd1902: TDATA = 50'b01100001110000000111101110100001110010001011011110;
        12'd1903: TDATA = 50'b01100001101111010101000110100001110001010110111111;
        12'd1904: TDATA = 50'b01100001101110100010011110100001110000100010100001;
        12'd1905: TDATA = 50'b01100001101101101111110110100001101111101110000011;
        12'd1906: TDATA = 50'b01100001101100111101001110100001101110111001100111;
        12'd1907: TDATA = 50'b01100001101100001010100110100001101110000101001100;
        12'd1908: TDATA = 50'b01100001101011011000000010100001101101010000110100;
        12'd1909: TDATA = 50'b01100001101010100101100000100001101100011100100000;
        12'd1910: TDATA = 50'b01100001101001110010111110100001101011101000001110;
        12'd1911: TDATA = 50'b01100001101001000000011100100001101010110011111100;
        12'd1912: TDATA = 50'b01100001101000001101111100100001101001111111101110;
        12'd1913: TDATA = 50'b01100001100111011011011110100001101001001011100001;
        12'd1914: TDATA = 50'b01100001100110101001000010100001101000010111011000;
        12'd1915: TDATA = 50'b01100001100101110110100110100001100111100011001111;
        12'd1916: TDATA = 50'b01100001100101000100001010100001100110101111001000;
        12'd1917: TDATA = 50'b01100001100100010001110100100001100101111011000111;
        12'd1918: TDATA = 50'b01100001100011011111011010100001100101000111000101;
        12'd1919: TDATA = 50'b01100001100010101101000010100001100100010011000011;
        12'd1920: TDATA = 50'b01100001100001111010101110100001100011011111001000;
        12'd1921: TDATA = 50'b01100001100001001000010110100001100010101011001000;
        12'd1922: TDATA = 50'b01100001100000010110000110100001100001110111010001;
        12'd1923: TDATA = 50'b01100001011111100011110010100001100001000011011001;
        12'd1924: TDATA = 50'b01100001011110110001100010100001100000001111100101;
        12'd1925: TDATA = 50'b01100001011101111111010010100001011111011011110001;
        12'd1926: TDATA = 50'b01100001011101001101000010100001011110100111111111;
        12'd1927: TDATA = 50'b01100001011100011010110110100001011101110100010000;
        12'd1928: TDATA = 50'b01100001011011101000101100100001011101000000100101;
        12'd1929: TDATA = 50'b01100001011010110110011110100001011100001100111000;
        12'd1930: TDATA = 50'b01100001011010000100011000100001011011011001010010;
        12'd1931: TDATA = 50'b01100001011001010010001010100001011010100101100110;
        12'd1932: TDATA = 50'b01100001011000100000000110100001011001110010000101;
        12'd1933: TDATA = 50'b01100001010111101110000000100001011000111110100001;
        12'd1934: TDATA = 50'b01100001010110111011111100100001011000001011000001;
        12'd1935: TDATA = 50'b01100001010110001001111000100001010111010111100010;
        12'd1936: TDATA = 50'b01100001010101010111110100100001010110100100000100;
        12'd1937: TDATA = 50'b01100001010100100101110010100001010101110000101010;
        12'd1938: TDATA = 50'b01100001010011110011110010100001010100111101010001;
        12'd1939: TDATA = 50'b01100001010011000001110100100001010100001001111011;
        12'd1940: TDATA = 50'b01100001010010001111110110100001010011010110100111;
        12'd1941: TDATA = 50'b01100001010001011101111010100001010010100011010110;
        12'd1942: TDATA = 50'b01100001010000101100000000100001010001110000000110;
        12'd1943: TDATA = 50'b01100001001111111010000100100001010000111100110111;
        12'd1944: TDATA = 50'b01100001001111001000001010100001010000001001101001;
        12'd1945: TDATA = 50'b01100001001110010110010100100001001111010110100010;
        12'd1946: TDATA = 50'b01100001001101100100100000100001001110100011011011;
        12'd1947: TDATA = 50'b01100001001100110010101010100001001101110000010110;
        12'd1948: TDATA = 50'b01100001001100000000110010100001001100111101001110;
        12'd1949: TDATA = 50'b01100001001011001111000100100001001100001010010000;
        12'd1950: TDATA = 50'b01100001001010011101001110100001001011010111001101;
        12'd1951: TDATA = 50'b01100001001001101011100000100001001010100100010000;
        12'd1952: TDATA = 50'b01100001001000111001110100100001001001110001011000;
        12'd1953: TDATA = 50'b01100001001000001000000010100001001000111110011011;
        12'd1954: TDATA = 50'b01100001000111010110010110100001001000001011100100;
        12'd1955: TDATA = 50'b01100001000110100100101010100001000111011000101110;
        12'd1956: TDATA = 50'b01100001000101110011000000100001000110100101111100;
        12'd1957: TDATA = 50'b01100001000101000001011000100001000101110011001011;
        12'd1958: TDATA = 50'b01100001000100001111101100100001000101000000010111;
        12'd1959: TDATA = 50'b01100001000011011110001000100001000100001101101110;
        12'd1960: TDATA = 50'b01100001000010101100100000100001000011011010111111;
        12'd1961: TDATA = 50'b01100001000001111011000000100001000010101000011010;
        12'd1962: TDATA = 50'b01100001000001001001011010100001000001110101110000;
        12'd1963: TDATA = 50'b01100001000000010111111010100001000001000011001101;
        12'd1964: TDATA = 50'b01100000111111100110010100100001000000010000100101;
        12'd1965: TDATA = 50'b01100000111110110100111010100000111111011110001001;
        12'd1966: TDATA = 50'b01100000111110000011011010100000111110101011101001;
        12'd1967: TDATA = 50'b01100000111101010001111010100000111101111001001001;
        12'd1968: TDATA = 50'b01100000111100100000011100100000111101000110101101;
        12'd1969: TDATA = 50'b01100000111011101111000110100000111100010100011000;
        12'd1970: TDATA = 50'b01100000111010111101101000100000111011100001111101;
        12'd1971: TDATA = 50'b01100000111010001100010010100000111010101111101010;
        12'd1972: TDATA = 50'b01100000111001011010111010100000111001111101010111;
        12'd1973: TDATA = 50'b01100000111000101001100100100000111001001011000101;
        12'd1974: TDATA = 50'b01100000110111111000001100100000111000011000110100;
        12'd1975: TDATA = 50'b01100000110111000110111000100000110111100110100111;
        12'd1976: TDATA = 50'b01100000110110010101101000100000110110110100011101;
        12'd1977: TDATA = 50'b01100000110101100100010110100000110110000010010101;
        12'd1978: TDATA = 50'b01100000110100110011000110100000110101010000001101;
        12'd1979: TDATA = 50'b01100000110100000001110100100000110100011110000110;
        12'd1980: TDATA = 50'b01100000110011010000100110100000110011101100000011;
        12'd1981: TDATA = 50'b01100000110010011111011100100000110010111010000011;
        12'd1982: TDATA = 50'b01100000110001101110001110100000110010001000000010;
        12'd1983: TDATA = 50'b01100000110000111101000010100000110001010110000100;
        12'd1984: TDATA = 50'b01100000110000001011111010100000110000100100001010;
        12'd1985: TDATA = 50'b01100000101111011010110010100000101111110010010001;
        12'd1986: TDATA = 50'b01100000101110101001101010100000101111000000011000;
        12'd1987: TDATA = 50'b01100000101101111000100110100000101110001110100100;
        12'd1988: TDATA = 50'b01100000101101000111100000100000101101011100110000;
        12'd1989: TDATA = 50'b01100000101100010110011110100000101100101011000000;
        12'd1990: TDATA = 50'b01100000101011100101011010100000101011111001001110;
        12'd1991: TDATA = 50'b01100000101010110100011000100000101011000111100000;
        12'd1992: TDATA = 50'b01100000101010000011011000100000101010010101110110;
        12'd1993: TDATA = 50'b01100000101001010010011010100000101001100100001100;
        12'd1994: TDATA = 50'b01100000101000100001011110100000101000110010100110;
        12'd1995: TDATA = 50'b01100000100111110000011110100000101000000000111110;
        12'd1996: TDATA = 50'b01100000100110111111100110100000100111001111011101;
        12'd1997: TDATA = 50'b01100000100110001110101010100000100110011101111001;
        12'd1998: TDATA = 50'b01100000100101011101110000100000100101101100011010;
        12'd1999: TDATA = 50'b01100000100100101100111010100000100100111010111110;
        12'd2000: TDATA = 50'b01100000100011111100000010100000100100001001100000;
        12'd2001: TDATA = 50'b01100000100011001011001110100000100011011000001000;
        12'd2002: TDATA = 50'b01100000100010011010010110100000100010100110101100;
        12'd2003: TDATA = 50'b01100000100001101001100110100000100001110101011001;
        12'd2004: TDATA = 50'b01100000100000111000110010100000100001000100000100;
        12'd2005: TDATA = 50'b01100000100000001000000010100000100000010010110011;
        12'd2006: TDATA = 50'b01100000011111010111010010100000011111100001100011;
        12'd2007: TDATA = 50'b01100000011110100110100010100000011110110000010011;
        12'd2008: TDATA = 50'b01100000011101110101110110100000011101111111001000;
        12'd2009: TDATA = 50'b01100000011101000101001100100000011101001110000000;
        12'd2010: TDATA = 50'b01100000011100010100011110100000011100011100110101;
        12'd2011: TDATA = 50'b01100000011011100011110010100000011011101011101100;
        12'd2012: TDATA = 50'b01100000011010110011001010100000011010111010101001;
        12'd2013: TDATA = 50'b01100000011010000010100100100000011010001001101000;
        12'd2014: TDATA = 50'b01100000011001010001111100100000011001011000100111;
        12'd2015: TDATA = 50'b01100000011000100001010110100000011000100111100110;
        12'd2016: TDATA = 50'b01100000010111110000110010100000010111110110101010;
        12'd2017: TDATA = 50'b01100000010111000000001110100000010111000101101110;
        12'd2018: TDATA = 50'b01100000010110001111101100100000010110010100110110;
        12'd2019: TDATA = 50'b01100000010101011111001100100000010101100011111111;
        12'd2020: TDATA = 50'b01100000010100101110101110100000010100110011001100;
        12'd2021: TDATA = 50'b01100000010011111110001100100000010100000010010110;
        12'd2022: TDATA = 50'b01100000010011001101101110100000010011010001100100;
        12'd2023: TDATA = 50'b01100000010010011101010100100000010010100000110110;
        12'd2024: TDATA = 50'b01100000010001101100111000100000010001110000001001;
        12'd2025: TDATA = 50'b01100000010000111100011110100000010000111111011101;
        12'd2026: TDATA = 50'b01100000010000001100000110100000010000001110110100;
        12'd2027: TDATA = 50'b01100000001111011011101110100000001111011110001100;
        12'd2028: TDATA = 50'b01100000001110101011010110100000001110101101100101;
        12'd2029: TDATA = 50'b01100000001101111011000100100000001101111101000100;
        12'd2030: TDATA = 50'b01100000001101001010101110100000001101001100100010;
        12'd2031: TDATA = 50'b01100000001100011010011010100000001100011100000000;
        12'd2032: TDATA = 50'b01100000001011101010001000100000001011101011100010;
        12'd2033: TDATA = 50'b01100000001010111001110110100000001010111011000100;
        12'd2034: TDATA = 50'b01100000001010001001100110100000001010001010101011;
        12'd2035: TDATA = 50'b01100000001001011001011000100000001001011010010010;
        12'd2036: TDATA = 50'b01100000001000101001001100100000001000101001111101;
        12'd2037: TDATA = 50'b01100000000111111001000000100000000111111001101000;
        12'd2038: TDATA = 50'b01100000000111001000110100100000000111001001010101;
        12'd2039: TDATA = 50'b01100000000110011000101000100000000110011001000010;
        12'd2040: TDATA = 50'b01100000000101101000011110100000000101101000110011;
        12'd2041: TDATA = 50'b01100000000100111000011000100000000100111000101000;
        12'd2042: TDATA = 50'b01100000000100001000010000100000000100001000011010;
        12'd2043: TDATA = 50'b01100000000011011000001100100000000011011000010100;
        12'd2044: TDATA = 50'b01100000000010101000000110100000000010101000001011;
        12'd2045: TDATA = 50'b01100000000001111000000100100000000001111000000101;
        12'd2046: TDATA = 50'b01100000000001001000000100100000000001001000000100;
        12'd2047: TDATA = 50'b01100000000000011000000000100000000000011000000000;
        12'd2048: TDATA = 50'b10111111111110100000000001111111111101000000000001;
        12'd2049: TDATA = 50'b10111111111011100000010001111111110111000000101011;
        12'd2050: TDATA = 50'b10111111111000100000011101111111110001000001011011;
        12'd2051: TDATA = 50'b10111111110101100000111011111111101011000010111011;
        12'd2052: TDATA = 50'b10111111110010100001011011111111100101000100101101;
        12'd2053: TDATA = 50'b10111111101111100010001001111111011111000111000011;
        12'd2054: TDATA = 50'b10111111101100100011000001111111011001001001111100;
        12'd2055: TDATA = 50'b10111111101001100100000001111111010011001101001101;
        12'd2056: TDATA = 50'b10111111100110100101000011111111001101010000110000;
        12'd2057: TDATA = 50'b10111111100011100110010111111111000111010101000011;
        12'd2058: TDATA = 50'b10111111100000100111110011111111000001011001110100;
        12'd2059: TDATA = 50'b10111111011101101001010011111110111011011110110110;
        12'd2060: TDATA = 50'b10111111011010101010111101111110110101100100010110;
        12'd2061: TDATA = 50'b10111111010111101100110001111110101111101010011010;
        12'd2062: TDATA = 50'b10111111010100101110101101111110101001110000110101;
        12'd2063: TDATA = 50'b10111111010001110000110011111110100011110111110011;
        12'd2064: TDATA = 50'b10111111001110110011000001111110011101111111001010;
        12'd2065: TDATA = 50'b10111111001011110101011001111110011000000111000100;
        12'd2066: TDATA = 50'b10111111001000110111111001111110010010001111010101;
        12'd2067: TDATA = 50'b10111111000101111010100011111110001100011000001010;
        12'd2068: TDATA = 50'b10111111000010111101010101111110000110100001010110;
        12'd2069: TDATA = 50'b10111111000000000000010001111110000000101011000101;
        12'd2070: TDATA = 50'b10111110111101000011010001111101111010110101000111;
        12'd2071: TDATA = 50'b10111110111010000110100001111101110100111111110001;
        12'd2072: TDATA = 50'b10111110110111001001111001111101101111001010111001;
        12'd2073: TDATA = 50'b10111110110100001101010001111101101001010110001100;
        12'd2074: TDATA = 50'b10111110110001010000110111111101100011100010001000;
        12'd2075: TDATA = 50'b10111110101110010100100101111101011101101110011100;
        12'd2076: TDATA = 50'b10111110101011011000100001111101010111111011011000;
        12'd2077: TDATA = 50'b10111110101000011100011101111101010010001000100000;
        12'd2078: TDATA = 50'b10111110100101100000101011111101001100010110011000;
        12'd2079: TDATA = 50'b10111110100010100100111011111101000110100100100000;
        12'd2080: TDATA = 50'b10111110011111101001010011111101000000110010111111;
        12'd2081: TDATA = 50'b10111110011100101101111001111100111011000010001000;
        12'd2082: TDATA = 50'b10111110011001110010100101111100110101010001100111;
        12'd2083: TDATA = 50'b10111110010110110111011001111100101111100001100100;
        12'd2084: TDATA = 50'b10111110010011111100010101111100101001110001110111;
        12'd2085: TDATA = 50'b10111110010001000001011011111100100100000010101110;
        12'd2086: TDATA = 50'b10111110001110000110101001111100011110010011111100;
        12'd2087: TDATA = 50'b10111110001011001100000001111100011000100101101100;
        12'd2088: TDATA = 50'b10111110001000010001011011111100010010110111101000;
        12'd2089: TDATA = 50'b10111110000101010111000011111100001101001010001100;
        12'd2090: TDATA = 50'b10111110000010011100111001111100000111011101011001;
        12'd2091: TDATA = 50'b10111101111111100010110011111100000001110000110110;
        12'd2092: TDATA = 50'b10111101111100101000110011111011111100000100101011;
        12'd2093: TDATA = 50'b10111101111001101110111001111011110110011000110111;
        12'd2094: TDATA = 50'b10111101110110110101001111111011110000101101101011;
        12'd2095: TDATA = 50'b10111101110011111011101001111011101011000010110110;
        12'd2096: TDATA = 50'b10111101110001000010010001111011100101011000100011;
        12'd2097: TDATA = 50'b10111101101110001000111011111011011111101110100010;
        12'd2098: TDATA = 50'b10111101101011001111101011111011011010000100110111;
        12'd2099: TDATA = 50'b10111101101000010110101101111011010100011011111010;
        12'd2100: TDATA = 50'b10111101100101011101110001111011001110110011001110;
        12'd2101: TDATA = 50'b10111101100010100100111111111011001001001010111111;
        12'd2102: TDATA = 50'b10111101011111101100010111111011000011100011001100;
        12'd2103: TDATA = 50'b10111101011100110011110111111010111101111011110101;
        12'd2104: TDATA = 50'b10111101011001111011011101111010111000010100110110;
        12'd2105: TDATA = 50'b10111101010111000011001111111010110010101110011000;
        12'd2106: TDATA = 50'b10111101010100001011000111111010101101001000010001;
        12'd2107: TDATA = 50'b10111101010001010011000101111010100111100010100001;
        12'd2108: TDATA = 50'b10111101001110011011001111111010100001111101010011;
        12'd2109: TDATA = 50'b10111101001011100011011111111010011100011000011011;
        12'd2110: TDATA = 50'b10111101001000101011111011111010010110110100000101;
        12'd2111: TDATA = 50'b10111101000101110100011101111010010001010000000110;
        12'd2112: TDATA = 50'b10111101000010111101000101111010001011101100011101;
        12'd2113: TDATA = 50'b10111101000000000101110011111010000110001001001011;
        12'd2114: TDATA = 50'b10111100111101001110101111111010000000100110100001;
        12'd2115: TDATA = 50'b10111100111010010111111001111001111011000100011000;
        12'd2116: TDATA = 50'b10111100110111100001000001111001110101100010011010;
        12'd2117: TDATA = 50'b10111100110100101010010011111001110000000000111000;
        12'd2118: TDATA = 50'b10111100110001110011101111111001101010011111110011;
        12'd2119: TDATA = 50'b10111100101110111101011001111001100100111111010101;
        12'd2120: TDATA = 50'b10111100101100000111000011111001011111011111000010;
        12'd2121: TDATA = 50'b10111100101001010000110011111001011001111111000100;
        12'd2122: TDATA = 50'b10111100100110011010110101111001010100011111110101;
        12'd2123: TDATA = 50'b10111100100011100100111001111001001111000000110101;
        12'd2124: TDATA = 50'b10111100100000101111000111111001001001100010010010;
        12'd2125: TDATA = 50'b10111100011101111001011111111001000100000100001010;
        12'd2126: TDATA = 50'b10111100011011000011111011111000111110100110011001;
        12'd2127: TDATA = 50'b10111100011000001110100001111000111001001001000011;
        12'd2128: TDATA = 50'b10111100010101011001010001111000110011101100001010;
        12'd2129: TDATA = 50'b10111100010010100100000011111000101110001111100000;
        12'd2130: TDATA = 50'b10111100001111101111000111111000101000110011100100;
        12'd2131: TDATA = 50'b10111100001100111010010001111000100011010111111101;
        12'd2132: TDATA = 50'b10111100001010000101011011111000011101111100100001;
        12'd2133: TDATA = 50'b10111100000111010000110001111000011000100001100111;
        12'd2134: TDATA = 50'b10111100000100011100001111111000010011000111001000;
        12'd2135: TDATA = 50'b10111100000001100111110111111000001101101101000101;
        12'd2136: TDATA = 50'b10111011111110110011100011111000001000010011010010;
        12'd2137: TDATA = 50'b10111011111011111111011101111000000010111010000110;
        12'd2138: TDATA = 50'b10111011111001001011011101110111111101100001010000;
        12'd2139: TDATA = 50'b10111011110110010111101001110111111000001000111011;
        12'd2140: TDATA = 50'b10111011110011100011110101110111110010110000110000;
        12'd2141: TDATA = 50'b10111011110000110000001111110111101101011001001101;
        12'd2142: TDATA = 50'b10111011101101111100110001110111101000000001111111;
        12'd2143: TDATA = 50'b10111011101011001001010101110111100010101011000001;
        12'd2144: TDATA = 50'b10111011101000010110000101110111011101010100100101;
        12'd2145: TDATA = 50'b10111011100101100010111011110111010111111110011110;
        12'd2146: TDATA = 50'b10111011100010101111111101110111010010101000111000;
        12'd2147: TDATA = 50'b10111011011111111101000101110111001101010011100111;
        12'd2148: TDATA = 50'b10111011011101001010010011110111000111111110101101;
        12'd2149: TDATA = 50'b10111011011010010111101101110111000010101010010011;
        12'd2150: TDATA = 50'b10111011010111100101001101110110111101010110001111;
        12'd2151: TDATA = 50'b10111011010100110010111001110110111000000010101100;
        12'd2152: TDATA = 50'b10111011010010000000100101110110110010101111010011;
        12'd2153: TDATA = 50'b10111011001111001110011101110110101101011100011011;
        12'd2154: TDATA = 50'b10111011001100011100100001110110101000001010000100;
        12'd2155: TDATA = 50'b10111011001001101010100101110110100010110111110111;
        12'd2156: TDATA = 50'b10111011000110111000110101110110011101100110001010;
        12'd2157: TDATA = 50'b10111011000100000111001011110110011000010100110100;
        12'd2158: TDATA = 50'b10111011000001010101101101110110010011000011111101;
        12'd2159: TDATA = 50'b10111010111110100100010101110110001101110011011101;
        12'd2160: TDATA = 50'b10111010111011110010111111110110001000100011001100;
        12'd2161: TDATA = 50'b10111010111001000001111001110110000011010011100001;
        12'd2162: TDATA = 50'b10111010110110010000111001110101111110000100001100;
        12'd2163: TDATA = 50'b10111010110011011111111101110101111000110101000110;
        12'd2164: TDATA = 50'b10111010110000101111001111110101110011100110100110;
        12'd2165: TDATA = 50'b10111010101101111110100011110101101110011000010111;
        12'd2166: TDATA = 50'b10111010101011001110000001110101101001001010100001;
        12'd2167: TDATA = 50'b10111010101000011101101001110101100011111101000111;
        12'd2168: TDATA = 50'b10111010100101101101011001110101011110110000001000;
        12'd2169: TDATA = 50'b10111010100010111101001111110101011001100011011110;
        12'd2170: TDATA = 50'b10111010100000001101000111110101010100010111000011;
        12'd2171: TDATA = 50'b10111010011101011101001111110101001111001011001111;
        12'd2172: TDATA = 50'b10111010011010101101011011110101001001111111101010;
        12'd2173: TDATA = 50'b10111010010111111101110001110101000100110100100101;
        12'd2174: TDATA = 50'b10111010010101001110001111110100111111101001110101;
        12'd2175: TDATA = 50'b10111010010010011110110101110100111010011111100000;
        12'd2176: TDATA = 50'b10111010001111101111100001110100110101010101100000;
        12'd2177: TDATA = 50'b10111010001101000000010011110100110000001011110101;
        12'd2178: TDATA = 50'b10111010001010010001010001110100101011000010101010;
        12'd2179: TDATA = 50'b10111010000111100010010001110100100101111001101111;
        12'd2180: TDATA = 50'b10111010000100110011011111110100100000110001010100;
        12'd2181: TDATA = 50'b10111010000010000100110001110100011011101001001101;
        12'd2182: TDATA = 50'b10111001111111010110001011110100010110100001011100;
        12'd2183: TDATA = 50'b10111001111100100111101101110100010001011010000101;
        12'd2184: TDATA = 50'b10111001111001111001010111110100001100010011001000;
        12'd2185: TDATA = 50'b10111001110111001011000011110100000111001100010110;
        12'd2186: TDATA = 50'b10111001110100011100111111110100000010000110001110;
        12'd2187: TDATA = 50'b10111001110001101110111111110011111101000000010101;
        12'd2188: TDATA = 50'b10111001101111000001001011110011110111111010111101;
        12'd2189: TDATA = 50'b10111001101100010011011011110011110010110101110100;
        12'd2190: TDATA = 50'b10111001101001100101110011110011101101110001000101;
        12'd2191: TDATA = 50'b10111001100110111000010001110011101000101100101010;
        12'd2192: TDATA = 50'b10111001100100001010110111110011100011101000101010;
        12'd2193: TDATA = 50'b10111001100001011101100101110011011110100100111111;
        12'd2194: TDATA = 50'b10111001011110110000011011110011011001100001101110;
        12'd2195: TDATA = 50'b10111001011100000011011001110011010100011110110111;
        12'd2196: TDATA = 50'b10111001011001010110011111110011001111011100010101;
        12'd2197: TDATA = 50'b10111001010110101001101001110011001010011010000111;
        12'd2198: TDATA = 50'b10111001010011111100111011110011000101011000001110;
        12'd2199: TDATA = 50'b10111001010001010000010111110011000000010110110101;
        12'd2200: TDATA = 50'b10111001001110100100000001110010111011010101111011;
        12'd2201: TDATA = 50'b10111001001011110111101001110010110110010101001010;
        12'd2202: TDATA = 50'b10111001001001001011011011110010110001010100110100;
        12'd2203: TDATA = 50'b10111001000110011111010111110010101100010100111000;
        12'd2204: TDATA = 50'b10111001000011110011010101110010100111010101001010;
        12'd2205: TDATA = 50'b10111001000001000111011111110010100010010101111101;
        12'd2206: TDATA = 50'b10111000111110011011101111110010011101010111000011;
        12'd2207: TDATA = 50'b10111000111011110000000101110010011000011000011110;
        12'd2208: TDATA = 50'b10111000111001000100100111110010010011011010011000;
        12'd2209: TDATA = 50'b10111000110110011001001111110010001110011100100111;
        12'd2210: TDATA = 50'b10111000110011101101111001110010001001011111000101;
        12'd2211: TDATA = 50'b10111000110001000010110001110010000100100010000010;
        12'd2212: TDATA = 50'b10111000101110010111100111110001111111100101001000;
        12'd2213: TDATA = 50'b10111000101011101100110011110001111010101000111110;
        12'd2214: TDATA = 50'b10111000101001000001111001110001110101101100110010;
        12'd2215: TDATA = 50'b10111000100110010111001111110001110000110001001011;
        12'd2216: TDATA = 50'b10111000100011101100101001110001101011110101111001;
        12'd2217: TDATA = 50'b10111000100001000010001011110001100110111010111010;
        12'd2218: TDATA = 50'b10111000011110010111110101110001100010000000010101;
        12'd2219: TDATA = 50'b10111000011011101101100101110001011101000110000101;
        12'd2220: TDATA = 50'b10111000011001000011011011110001011000001100001000;
        12'd2221: TDATA = 50'b10111000010110011001011101110001010011010010101011;
        12'd2222: TDATA = 50'b10111000010011101111100001110001001110011001011100;
        12'd2223: TDATA = 50'b10111000010001000101110011110001001001100000101100;
        12'd2224: TDATA = 50'b10111000001110011100000111110001000100101000001011;
        12'd2225: TDATA = 50'b10111000001011110010100111110000111111110000001001;
        12'd2226: TDATA = 50'b10111000001001001001001001110000111010111000010101;
        12'd2227: TDATA = 50'b10111000000110011111110011110000110110000000110110;
        12'd2228: TDATA = 50'b10111000000011110110100101110000110001001001110000;
        12'd2229: TDATA = 50'b10111000000001001101011111110000101100010011000011;
        12'd2230: TDATA = 50'b10110111111110100100100011110000100111011100110000;
        12'd2231: TDATA = 50'b10110111111011111011101011110000100010100110101011;
        12'd2232: TDATA = 50'b10110111111001010010111011110000011101110001000000;
        12'd2233: TDATA = 50'b10110111110110101010010001110000011000111011101000;
        12'd2234: TDATA = 50'b10110111110100000001101111110000010100000110101010;
        12'd2235: TDATA = 50'b10110111110001011001010101110000001111010010000000;
        12'd2236: TDATA = 50'b10110111101110110000111111110000001010011101101010;
        12'd2237: TDATA = 50'b10110111101100001000111001110000000101101001110111;
        12'd2238: TDATA = 50'b10110111101001100000110011110000000000110110001110;
        12'd2239: TDATA = 50'b10110111100110111000110011101111111100000010111000;
        12'd2240: TDATA = 50'b10110111100100010000111001101111110111001111110111;
        12'd2241: TDATA = 50'b10110111100001101001001011101111110010011101010100;
        12'd2242: TDATA = 50'b10110111011111000001100011101111101101101011000100;
        12'd2243: TDATA = 50'b10110111011100011010000001101111101000111001001000;
        12'd2244: TDATA = 50'b10110111011001110010101001101111100100000111100110;
        12'd2245: TDATA = 50'b10110111010111001011011001101111011111010110011100;
        12'd2246: TDATA = 50'b10110111010100100100001111101111011010100101100111;
        12'd2247: TDATA = 50'b10110111010001111101000101101111010101110100111001;
        12'd2248: TDATA = 50'b10110111001111010110001001101111010001000100110000;
        12'd2249: TDATA = 50'b10110111001100101111010101101111001100010100111011;
        12'd2250: TDATA = 50'b10110111001010001000100011101111000111100101010011;
        12'd2251: TDATA = 50'b10110111000111100001111101101111000010110110001010;
        12'd2252: TDATA = 50'b10110111000100111011011101101110111110000111010101;
        12'd2253: TDATA = 50'b10110111000010010101000011101110111001011000110011;
        12'd2254: TDATA = 50'b10110110111111101110110001101110110100101010101010;
        12'd2255: TDATA = 50'b10110110111101001000100111101110101111111100110101;
        12'd2256: TDATA = 50'b10110110111010100010100001101110101011001111010011;
        12'd2257: TDATA = 50'b10110110110111111100101001101110100110100010001111;
        12'd2258: TDATA = 50'b10110110110101010110101101101110100001110101001110;
        12'd2259: TDATA = 50'b10110110110010110000111111101110011101001000110001;
        12'd2260: TDATA = 50'b10110110110000001011010011101110011000011100011101;
        12'd2261: TDATA = 50'b10110110101101100101110101101110010011110000101100;
        12'd2262: TDATA = 50'b10110110101011000000011101101110001111000101001111;
        12'd2263: TDATA = 50'b10110110101000011011000111101110001010011001111111;
        12'd2264: TDATA = 50'b10110110100101110101111111101110000101101111001110;
        12'd2265: TDATA = 50'b10110110100011010000111011101110000001000100110000;
        12'd2266: TDATA = 50'b10110110100000101011111011101101111100011010100000;
        12'd2267: TDATA = 50'b10110110011110000111000001101101110111110000100011;
        12'd2268: TDATA = 50'b10110110011011100010010011101101110011000111000100;
        12'd2269: TDATA = 50'b10110110011000111101101001101101101110011101110011;
        12'd2270: TDATA = 50'b10110110010110011001000011101101101001110100110101;
        12'd2271: TDATA = 50'b10110110010011110100101011101101100101001100010110;
        12'd2272: TDATA = 50'b10110110010001010000010101101101100000100100000100;
        12'd2273: TDATA = 50'b10110110001110101100000111101101011011111100001010;
        12'd2274: TDATA = 50'b10110110001100001000000001101101010111010100100100;
        12'd2275: TDATA = 50'b10110110001001100011111111101101010010101101010001;
        12'd2276: TDATA = 50'b10110110000111000000001011101101001110000110011011;
        12'd2277: TDATA = 50'b10110110000100011100011001101101001001011111110100;
        12'd2278: TDATA = 50'b10110110000001111000101101101101000100111001011111;
        12'd2279: TDATA = 50'b10110101111111010101001001101101000000010011100011;
        12'd2280: TDATA = 50'b10110101111100110001101101101100111011101101111010;
        12'd2281: TDATA = 50'b10110101111010001110011001101100110111001000101001;
        12'd2282: TDATA = 50'b10110101110111101011000101101100110010100011100001;
        12'd2283: TDATA = 50'b10110101110101000111111101101100101101111110110110;
        12'd2284: TDATA = 50'b10110101110010100101000001101100101001011010101001;
        12'd2285: TDATA = 50'b10110101110000000010000001101100100100110110011111;
        12'd2286: TDATA = 50'b10110101101101011111001111101100100000010010110010;
        12'd2287: TDATA = 50'b10110101101010111100100001101100011011101111011001;
        12'd2288: TDATA = 50'b10110101101000011001111011101100010111001100010010;
        12'd2289: TDATA = 50'b10110101100101110111011101101100010010101001100011;
        12'd2290: TDATA = 50'b10110101100011010101000101101100001110000111001000;
        12'd2291: TDATA = 50'b10110101100000110010101111101100001001100100111010;
        12'd2292: TDATA = 50'b10110101011110010000101001101100000101000011001110;
        12'd2293: TDATA = 50'b10110101011011101110100011101100000000100001101011;
        12'd2294: TDATA = 50'b10110101011001001100100111101011111100000000100000;
        12'd2295: TDATA = 50'b10110101010110101010101001101011110111011111011101;
        12'd2296: TDATA = 50'b10110101010100001000111111101011110010111111000011;
        12'd2297: TDATA = 50'b10110101010001100111010011101011101110011110110000;
        12'd2298: TDATA = 50'b10110101001111000101110001101011101001111110110101;
        12'd2299: TDATA = 50'b10110101001100100100011001101011100101011111010011;
        12'd2300: TDATA = 50'b10110101001010000011000011101011100000111111111101;
        12'd2301: TDATA = 50'b10110101000111100001110011101011011100100000111011;
        12'd2302: TDATA = 50'b10110101000101000000101111101011011000000010010110;
        12'd2303: TDATA = 50'b10110101000010011111110001101011010011100100000011;
        12'd2304: TDATA = 50'b10110100111111111110110011101011001111000101111000;
        12'd2305: TDATA = 50'b10110100111101011101111011101011001010101000000000;
        12'd2306: TDATA = 50'b10110100111010111101010001101011000110001010101011;
        12'd2307: TDATA = 50'b10110100111000011100101111101011000001101101101000;
        12'd2308: TDATA = 50'b10110100110101111100001111101010111101010000110010;
        12'd2309: TDATA = 50'b10110100110011011011110101101010111000110100001111;
        12'd2310: TDATA = 50'b10110100110000111011100011101010110100011000000100;
        12'd2311: TDATA = 50'b10110100101110011011011001101010101111111100001011;
        12'd2312: TDATA = 50'b10110100101011111011010011101010101011100000100101;
        12'd2313: TDATA = 50'b10110100101001011011010101101010100111000101010001;
        12'd2314: TDATA = 50'b10110100100110111011011111101010100010101010010101;
        12'd2315: TDATA = 50'b10110100100100011011101111101010011110001111101011;
        12'd2316: TDATA = 50'b10110100100001111100000001101010011001110101001110;
        12'd2317: TDATA = 50'b10110100011111011100100001101010010101011011001111;
        12'd2318: TDATA = 50'b10110100011100111101000011101010010001000001011101;
        12'd2319: TDATA = 50'b10110100011010011101101011101010001100100111111100;
        12'd2320: TDATA = 50'b10110100010111111110100001101010001000001110111111;
        12'd2321: TDATA = 50'b10110100010101011111001111101010000011110101111001;
        12'd2322: TDATA = 50'b10110100010011000000001111101001111111011101011010;
        12'd2323: TDATA = 50'b10110100010000100001011001101001111011000101010100;
        12'd2324: TDATA = 50'b10110100001110000010100001101001110110101101010100;
        12'd2325: TDATA = 50'b10110100001011100011110011101001110010010101101101;
        12'd2326: TDATA = 50'b10110100001001000101001001101001101101111110010010;
        12'd2327: TDATA = 50'b10110100000110100110100111101001101001100111001111;
        12'd2328: TDATA = 50'b10110100000100001000001011101001100101010000011110;
        12'd2329: TDATA = 50'b10110100000001101001110111101001100000111010000101;
        12'd2330: TDATA = 50'b10110011111111001011101011101001011100100011111110;
        12'd2331: TDATA = 50'b10110011111100101101100001101001011000001110000100;
        12'd2332: TDATA = 50'b10110011111010001111011111101001010011111000100001;
        12'd2333: TDATA = 50'b10110011110111110001100101101001001111100011010000;
        12'd2334: TDATA = 50'b10110011110101010011110011101001001011001110010111;
        12'd2335: TDATA = 50'b10110011110010110110000111101001000110111001110000;
        12'd2336: TDATA = 50'b10110011110000011000011011101001000010100101010000;
        12'd2337: TDATA = 50'b10110011101101111011000001101000111110010001011000;
        12'd2338: TDATA = 50'b10110011101011011101100011101000111001111101100010;
        12'd2339: TDATA = 50'b10110011101001000000001101101000110101101001111110;
        12'd2340: TDATA = 50'b10110011100110100011000001101000110001010110110110;
        12'd2341: TDATA = 50'b10110011100100000101111001101000101101000011111011;
        12'd2342: TDATA = 50'b10110011100001101000111011101000101000110001011000;
        12'd2343: TDATA = 50'b10110011011111001011111111101000100100011111000001;
        12'd2344: TDATA = 50'b10110011011100101111001111101000100000001101000111;
        12'd2345: TDATA = 50'b10110011011010010010100001101000011011111011011001;
        12'd2346: TDATA = 50'b10110011010111110101111011101000010111101001111101;
        12'd2347: TDATA = 50'b10110011010101011001011101101000010011011000111001;
        12'd2348: TDATA = 50'b10110011010010111101000001101000001111001000000001;
        12'd2349: TDATA = 50'b10110011010000100000101101101000001010110111011011;
        12'd2350: TDATA = 50'b10110011001110000100011011101000000110100111000010;
        12'd2351: TDATA = 50'b10110011001011101000010111101000000010010111001010;
        12'd2352: TDATA = 50'b10110011001001001100010101100111111110000111011010;
        12'd2353: TDATA = 50'b10110011000110110000100001100111111001111000001011;
        12'd2354: TDATA = 50'b10110011000100010100101001100111110101101000111110;
        12'd2355: TDATA = 50'b10110011000001111000111011100111110001011010001001;
        12'd2356: TDATA = 50'b10110010111111011101010011100111101101001011100101;
        12'd2357: TDATA = 50'b10110010111101000001110111100111101000111101011101;
        12'd2358: TDATA = 50'b10110010111010100110011001100111100100101111011000;
        12'd2359: TDATA = 50'b10110010111000001011001001100111100000100001110011;
        12'd2360: TDATA = 50'b10110010110101101111111001100111011100010100010111;
        12'd2361: TDATA = 50'b10110010110011010100110001100111011000000111010001;
        12'd2362: TDATA = 50'b10110010110000111001110001100111010011111010011100;
        12'd2363: TDATA = 50'b10110010101110011110111001100111001111101101111111;
        12'd2364: TDATA = 50'b10110010101100000100000001100111001011100001101001;
        12'd2365: TDATA = 50'b10110010101001101001010001100111000111010101101010;
        12'd2366: TDATA = 50'b10110010100111001110101011100111000011001010000001;
        12'd2367: TDATA = 50'b10110010100100110100001011100110111110111110101010;
        12'd2368: TDATA = 50'b10110010100010011001110001100110111010110011100101;
        12'd2369: TDATA = 50'b10110010011111111111010111100110110110101000100111;
        12'd2370: TDATA = 50'b10110010011101100101001001100110110010011110000101;
        12'd2371: TDATA = 50'b10110010011011001011000001100110101110010011110101;
        12'd2372: TDATA = 50'b10110010011000110000111111100110101010001001110110;
        12'd2373: TDATA = 50'b10110010010110010111000011100110100110000000001001;
        12'd2374: TDATA = 50'b10110010010011111101010001100110100001110110110010;
        12'd2375: TDATA = 50'b10110010010001100011100001100110011101101101100111;
        12'd2376: TDATA = 50'b10110010001111001001110011100110011001100100101001;
        12'd2377: TDATA = 50'b10110010001100110000010011100110010101011100000111;
        12'd2378: TDATA = 50'b10110010001010010110110101100110010001010011110001;
        12'd2379: TDATA = 50'b10110010000111111101011101100110001101001011101101;
        12'd2380: TDATA = 50'b10110010000101100100001011100110001001000011111010;
        12'd2381: TDATA = 50'b10110010000011001011000001100110000100111100011101;
        12'd2382: TDATA = 50'b10110010000000110001111111100110000000110101010010;
        12'd2383: TDATA = 50'b10110001111110011000111111100101111100101110010011;
        12'd2384: TDATA = 50'b10110001111100000000000101100101111000100111100101;
        12'd2385: TDATA = 50'b10110001111001100111010111100101110100100001010100;
        12'd2386: TDATA = 50'b10110001110111001110101011100101110000011011001110;
        12'd2387: TDATA = 50'b10110001110100110110000011100101101100010101010100;
        12'd2388: TDATA = 50'b10110001110010011101100111100101101000001111110111;
        12'd2389: TDATA = 50'b10110001110000000101001011100101100100001010100000;
        12'd2390: TDATA = 50'b10110001101101101100111001100101100000000101011111;
        12'd2391: TDATA = 50'b10110001101011010100101011100101011100000000110000;
        12'd2392: TDATA = 50'b10110001101000111100100101100101010111111100010010;
        12'd2393: TDATA = 50'b10110001100110100100100011100101010011111000000101;
        12'd2394: TDATA = 50'b10110001100100001100101011100101001111110100001111;
        12'd2395: TDATA = 50'b10110001100001110100110111100101001011110000100101;
        12'd2396: TDATA = 50'b10110001011111011101000111100101000111101101001011;
        12'd2397: TDATA = 50'b10110001011101000101011111100101000011101010000100;
        12'd2398: TDATA = 50'b10110001011010101101111011100100111111100111001101;
        12'd2399: TDATA = 50'b10110001011000010110011111100100111011100100100111;
        12'd2400: TDATA = 50'b10110001010101111111000111100100110111100010010011;
        12'd2401: TDATA = 50'b10110001010011100111111001100100110011100000010100;
        12'd2402: TDATA = 50'b10110001010001010000101111100100101111011110100010;
        12'd2403: TDATA = 50'b10110001001110111001101001100100101011011101000001;
        12'd2404: TDATA = 50'b10110001001100100010101011100100100111011011110001;
        12'd2405: TDATA = 50'b10110001001010001011110101100100100011011010110111;
        12'd2406: TDATA = 50'b10110001000111110100111111100100011111011010000100;
        12'd2407: TDATA = 50'b10110001000101011110010101100100011011011001101100;
        12'd2408: TDATA = 50'b10110001000011000111101011100100010111011001011011;
        12'd2409: TDATA = 50'b10110001000000110001001111100100010011011001101010;
        12'd2410: TDATA = 50'b10110000111110011010110101100100001111011010000000;
        12'd2411: TDATA = 50'b10110000111100000100011111100100001011011010101000;
        12'd2412: TDATA = 50'b10110000111001101110010111100100000111011011101010;
        12'd2413: TDATA = 50'b10110000110111011000000111100100000011011100101001;
        12'd2414: TDATA = 50'b10110000110101000010000111100011111111011110001000;
        12'd2415: TDATA = 50'b10110000110010101100001011100011111011011111110010;
        12'd2416: TDATA = 50'b10110000110000010110010111100011110111100001110011;
        12'd2417: TDATA = 50'b10110000101110000000101001100011110011100100000101;
        12'd2418: TDATA = 50'b10110000101011101011000001100011101111100110101000;
        12'd2419: TDATA = 50'b10110000101001010101011001100011101011101001010001;
        12'd2420: TDATA = 50'b10110000100110111111111001100011100111101100010000;
        12'd2421: TDATA = 50'b10110000100100101010100001100011100011101111100000;
        12'd2422: TDATA = 50'b10110000100010010101001011100011011111110010111100;
        12'd2423: TDATA = 50'b10110000011111111111111011100011011011110110101001;
        12'd2424: TDATA = 50'b10110000011101101010111001100011010111111010110110;
        12'd2425: TDATA = 50'b10110000011011010101111001100011010011111111001001;
        12'd2426: TDATA = 50'b10110000011001000000111011100011010000000011101000;
        12'd2427: TDATA = 50'b10110000010110101100001001100011001100001000100010;
        12'd2428: TDATA = 50'b10110000010100010111011001100011001000001101100111;
        12'd2429: TDATA = 50'b10110000010010000010110011100011000100010011000011;
        12'd2430: TDATA = 50'b10110000001111101110001011100011000000011000100000;
        12'd2431: TDATA = 50'b10110000001101011001110001100010111100011110011100;
        12'd2432: TDATA = 50'b10110000001011000101011001100010111000100100100101;
        12'd2433: TDATA = 50'b10110000001000110001001001100010110100101010111110;
        12'd2434: TDATA = 50'b10110000000110011100110111100010110000110001011110;
        12'd2435: TDATA = 50'b10110000000100001000110011100010101100111000011000;
        12'd2436: TDATA = 50'b10110000000001110100110011100010101000111111100011;
        12'd2437: TDATA = 50'b10101111111111100000110101100010100101000110110101;
        12'd2438: TDATA = 50'b10101111111101001101000101100010100001001110100110;
        12'd2439: TDATA = 50'b10101111111010111001010001100010011101010110011001;
        12'd2440: TDATA = 50'b10101111111000100101101011100010011001011110100110;
        12'd2441: TDATA = 50'b10101111110110010010000111100010010101100110111111;
        12'd2442: TDATA = 50'b10101111110011111110101001100010010001101111101001;
        12'd2443: TDATA = 50'b10101111110001101011010001100010001101111000100011;
        12'd2444: TDATA = 50'b10101111101111011000000001100010001010000001110010;
        12'd2445: TDATA = 50'b10101111101101000100101111100010000110001011000011;
        12'd2446: TDATA = 50'b10101111101010110001101101100010000010010100110100;
        12'd2447: TDATA = 50'b10101111101000011110101101100001111110011110110000;
        12'd2448: TDATA = 50'b10101111100110001011101111100001111010101000111000;
        12'd2449: TDATA = 50'b10101111100011111000111111100001110110110011011010;
        12'd2450: TDATA = 50'b10101111100001100110010001100001110010111110000111;
        12'd2451: TDATA = 50'b10101111011111010011101001100001101111001001000101;
        12'd2452: TDATA = 50'b10101111011101000001000001100001101011010100001001;
        12'd2453: TDATA = 50'b10101111011010101110100001100001100111011111100011;
        12'd2454: TDATA = 50'b10101111011000011100001001100001100011101011001101;
        12'd2455: TDATA = 50'b10101111010110001001111001100001011111110111001100;
        12'd2456: TDATA = 50'b10101111010011110111101011100001011100000011010111;
        12'd2457: TDATA = 50'b10101111010001100101100001100001011000001111101101;
        12'd2458: TDATA = 50'b10101111001111010011100001100001010100011100011001;
        12'd2459: TDATA = 50'b10101111001101000001101001100001010000101001011010;
        12'd2460: TDATA = 50'b10101111001010101111110001100001001100110110100001;
        12'd2461: TDATA = 50'b10101111001000011101111111100001001001000011111001;
        12'd2462: TDATA = 50'b10101111000110001100010011100001000101010001100000;
        12'd2463: TDATA = 50'b10101111000011111010101101100001000001011111011000;
        12'd2464: TDATA = 50'b10101111000001101001001101100000111101101101100001;
        12'd2465: TDATA = 50'b10101110111111010111111001100000111001111100000011;
        12'd2466: TDATA = 50'b10101110111101000110100001100000110110001010100111;
        12'd2467: TDATA = 50'b10101110111010110101010011100000110010011001100000;
        12'd2468: TDATA = 50'b10101110111000100100001011100000101110101000101001;
        12'd2469: TDATA = 50'b10101110110110010011000111100000101010110111111110;
        12'd2470: TDATA = 50'b10101110110100000010001011100000100111000111100111;
        12'd2471: TDATA = 50'b10101110110001110001010001100000100011010111011100;
        12'd2472: TDATA = 50'b10101110101111100000011111100000011111100111100001;
        12'd2473: TDATA = 50'b10101110101101001111110001100000011011110111110110;
        12'd2474: TDATA = 50'b10101110101010111111001011100000011000001000011011;
        12'd2475: TDATA = 50'b10101110101000101110101101100000010100011001010110;
        12'd2476: TDATA = 50'b10101110100110011110010001100000010000101010011011;
        12'd2477: TDATA = 50'b10101110100100001101111001100000001100111011101100;
        12'd2478: TDATA = 50'b10101110100001111101100111100000001001001101001101;
        12'd2479: TDATA = 50'b10101110011111101101100001100000000101011111000111;
        12'd2480: TDATA = 50'b10101110011101011101011011100000000001110001001000;
        12'd2481: TDATA = 50'b10101110011011001101011011011111111110000011011001;
        12'd2482: TDATA = 50'b10101110011000111101011111011111111010010101110101;
        12'd2483: TDATA = 50'b10101110010110101101100111011111110110101000100001;
        12'd2484: TDATA = 50'b10101110010100011101111001011111110010111011100010;
        12'd2485: TDATA = 50'b10101110010010001110001111011111101111001110101110;
        12'd2486: TDATA = 50'b10101110001111111110101101011111101011100010001111;
        12'd2487: TDATA = 50'b10101110001101101111010001011111100111110110000000;
        12'd2488: TDATA = 50'b10101110001011011111110101011111100100001001110110;
        12'd2489: TDATA = 50'b10101110001001010000100001011111100000011110000010;
        12'd2490: TDATA = 50'b10101110000111000001010101011111011100110010011110;
        12'd2491: TDATA = 50'b10101110000100110010001011011111011001000111000101;
        12'd2492: TDATA = 50'b10101110000010100011001001011111010101011100000000;
        12'd2493: TDATA = 50'b10101110000000010100001011011111010001110001000111;
        12'd2494: TDATA = 50'b10101101111110000101010011011111001110000110011101;
        12'd2495: TDATA = 50'b10101101111011110110100001011111001010011100000100;
        12'd2496: TDATA = 50'b10101101111001100111110011011111000110110001110101;
        12'd2497: TDATA = 50'b10101101110111011001001101011111000011000111111011;
        12'd2498: TDATA = 50'b10101101110101001010101101011110111111011110010001;
        12'd2499: TDATA = 50'b10101101110010111100001101011110111011110100101101;
        12'd2500: TDATA = 50'b10101101110000101101111001011110111000001011100010;
        12'd2501: TDATA = 50'b10101101101110011111100101011110110100100010011101;
        12'd2502: TDATA = 50'b10101101101100010001011001011110110000111001101101;
        12'd2503: TDATA = 50'b10101101101010000011010001011110101101010001001000;
        12'd2504: TDATA = 50'b10101101100111110101001111011110101001101000110011;
        12'd2505: TDATA = 50'b10101101100101100111010111011110100110000000110011;
        12'd2506: TDATA = 50'b10101101100011011001100001011110100010011000111101;
        12'd2507: TDATA = 50'b10101101100001001011110001011110011110110001010111;
        12'd2508: TDATA = 50'b10101101011110111110000001011110011011001001110111;
        12'd2509: TDATA = 50'b10101101011100110000011101011110010111100010110000;
        12'd2510: TDATA = 50'b10101101011010100010111011011110010011111011110100;
        12'd2511: TDATA = 50'b10101101011000010101100001011110010000010101001000;
        12'd2512: TDATA = 50'b10101101010110001000001011011110001100101110101011;
        12'd2513: TDATA = 50'b10101101010011111010111001011110001001001000011010;
        12'd2514: TDATA = 50'b10101101010001101101101011011110000101100010010010;
        12'd2515: TDATA = 50'b10101101001111100000100111011110000001111100100101;
        12'd2516: TDATA = 50'b10101101001101010011100111011101111110010111000010;
        12'd2517: TDATA = 50'b10101101001011000110110011011101111010110001111000;
        12'd2518: TDATA = 50'b10101101001000111001111001011101110111001100101011;
        12'd2519: TDATA = 50'b10101101000110101101001011011101110011100111110111;
        12'd2520: TDATA = 50'b10101101000100100000100001011101110000000011001101;
        12'd2521: TDATA = 50'b10101101000010010011111001011101101100011110101111;
        12'd2522: TDATA = 50'b10101101000000000111011001011101101000111010100100;
        12'd2523: TDATA = 50'b10101100111101111011000001011101100101010110101001;
        12'd2524: TDATA = 50'b10101100111011101110101011011101100001110010111001;
        12'd2525: TDATA = 50'b10101100111001100010011011011101011110001111011001;
        12'd2526: TDATA = 50'b10101100110111010110001011011101011010101011111110;
        12'd2527: TDATA = 50'b10101100110101001010001001011101010111001001000001;
        12'd2528: TDATA = 50'b10101100110010111110001001011101010011100110001010;
        12'd2529: TDATA = 50'b10101100110000110010010001011101010000000011100111;
        12'd2530: TDATA = 50'b10101100101110100110011001011101001100100001001010;
        12'd2531: TDATA = 50'b10101100101100011010101001011101001000111111000001;
        12'd2532: TDATA = 50'b10101100101010001110111011011101000101011100111110;
        12'd2533: TDATA = 50'b10101100101000000011010111011101000001111011010100;
        12'd2534: TDATA = 50'b10101100100101110111110111011100111110011001110101;
        12'd2535: TDATA = 50'b10101100100011101100100001011100111010111000101010;
        12'd2536: TDATA = 50'b10101100100001100001001001011100110111010111100100;
        12'd2537: TDATA = 50'b10101100011111010101111001011100110011110110101110;
        12'd2538: TDATA = 50'b10101100011101001010101011011100110000010110000011;
        12'd2539: TDATA = 50'b10101100011010111111100011011100101100110101100110;
        12'd2540: TDATA = 50'b10101100011000110100100111011100101001010101100011;
        12'd2541: TDATA = 50'b10101100010110101001101011011100100101110101100110;
        12'd2542: TDATA = 50'b10101100010100011110110101011100100010010101110111;
        12'd2543: TDATA = 50'b10101100010010010100000001011100011110110110010100;
        12'd2544: TDATA = 50'b10101100010000001001010111011100011011010111000100;
        12'd2545: TDATA = 50'b10101100001101111110110001011100010111110111111111;
        12'd2546: TDATA = 50'b10101100001011110100001111011100010100011001001001;
        12'd2547: TDATA = 50'b10101100001001101001110101011100010000111010100010;
        12'd2548: TDATA = 50'b10101100000111011111011101011100001101011100000101;
        12'd2549: TDATA = 50'b10101100000101010101000111011100001001111101110100;
        12'd2550: TDATA = 50'b10101100000011001011000001011100000110011111111111;
        12'd2551: TDATA = 50'b10101100000001000000111011011100000011000010010001;
        12'd2552: TDATA = 50'b10101011111110110110111011011011111111100100110001;
        12'd2553: TDATA = 50'b10101011111100101100111011011011111100000111010111;
        12'd2554: TDATA = 50'b10101011111010100011000001011011111000101010001100;
        12'd2555: TDATA = 50'b10101011111000011001010001011011110101001101010110;
        12'd2556: TDATA = 50'b10101011110110001111100011011011110001110000101001;
        12'd2557: TDATA = 50'b10101011110100000101111011011011101110010100001100;
        12'd2558: TDATA = 50'b10101011110001111100011001011011101010110111111110;
        12'd2559: TDATA = 50'b10101011101111110010111001011011100111011011111010;
        12'd2560: TDATA = 50'b10101011101101101001100001011011100100000000000101;
        12'd2561: TDATA = 50'b10101011101011100000001011011011100000100100011010;
        12'd2562: TDATA = 50'b10101011101001010110111011011011011101001000111111;
        12'd2563: TDATA = 50'b10101011100111001101110111011011011001101101111100;
        12'd2564: TDATA = 50'b10101011100101000100101111011011010110010010111010;
        12'd2565: TDATA = 50'b10101011100010111011110001011011010010111000001100;
        12'd2566: TDATA = 50'b10101011100000110010111001011011001111011101101101;
        12'd2567: TDATA = 50'b10101011011110101010000101011011001100000011011000;
        12'd2568: TDATA = 50'b10101011011100100001010011011011001000101001001101;
        12'd2569: TDATA = 50'b10101011011010011000101001011011000101001111010110;
        12'd2570: TDATA = 50'b10101011011000010000000111011011000001110101101110;
        12'd2571: TDATA = 50'b10101011010110000111100111011010111110011100010000;
        12'd2572: TDATA = 50'b10101011010011111111001001011010111011000010111100;
        12'd2573: TDATA = 50'b10101011010001110110110011011010110111101001111000;
        12'd2574: TDATA = 50'b10101011001111101110100001011010110100010001000010;
        12'd2575: TDATA = 50'b10101011001101100110011001011010110000111000100000;
        12'd2576: TDATA = 50'b10101011001011011110010001011010101101100000000011;
        12'd2577: TDATA = 50'b10101011001001010110001101011010101010000111110001;
        12'd2578: TDATA = 50'b10101011000111001110010011011010100110101111110111;
        12'd2579: TDATA = 50'b10101011000101000110100001011010100011011000001100;
        12'd2580: TDATA = 50'b10101011000010111110101011011010100000000000100001;
        12'd2581: TDATA = 50'b10101011000000110110111011011010011100101001000101;
        12'd2582: TDATA = 50'b10101010111110101111010001011010011001010001111001;
        12'd2583: TDATA = 50'b10101010111100100111101111011010010101111010111111;
        12'd2584: TDATA = 50'b10101010111010100000010001011010010010100100010000;
        12'd2585: TDATA = 50'b10101010111000011000111001011010001111001101110000;
        12'd2586: TDATA = 50'b10101010110110010001100001011010001011110111010101;
        12'd2587: TDATA = 50'b10101010110100001010001111011010001000100001001001;
        12'd2588: TDATA = 50'b10101010110010000011001001011010000101001011010101;
        12'd2589: TDATA = 50'b10101010101111111100000111011010000001110101101011;
        12'd2590: TDATA = 50'b10101010101101110101000011011001111110100000000110;
        12'd2591: TDATA = 50'b10101010101011101110000111011001111011001010110000;
        12'd2592: TDATA = 50'b10101010101001100111001111011001110111110101101001;
        12'd2593: TDATA = 50'b10101010100111100000100001011001110100100000110110;
        12'd2594: TDATA = 50'b10101010100101011001110011011001110001001100000111;
        12'd2595: TDATA = 50'b10101010100011010011001011011001101101110111101000;
        12'd2596: TDATA = 50'b10101010100001001100101001011001101010100011010111;
        12'd2597: TDATA = 50'b10101010011111000110010001011001100111001111011001;
        12'd2598: TDATA = 50'b10101010011100111111110101011001100011111011011100;
        12'd2599: TDATA = 50'b10101010011010111001100001011001100000100111110010;
        12'd2600: TDATA = 50'b10101010011000110011010101011001011101010100010111;
        12'd2601: TDATA = 50'b10101010010110101101001011011001011010000001000110;
        12'd2602: TDATA = 50'b10101010010100100111000111011001010110101110000100;
        12'd2603: TDATA = 50'b10101010010010100001001001011001010011011011010000;
        12'd2604: TDATA = 50'b10101010010000011011001011011001010000001000100010;
        12'd2605: TDATA = 50'b10101010001110010101010011011001001100110110000010;
        12'd2606: TDATA = 50'b10101010001100001111100111011001001001100011111010;
        12'd2607: TDATA = 50'b10101010001010001001111011011001000110010001110111;
        12'd2608: TDATA = 50'b10101010001000000100010001011001000010111111111110;
        12'd2609: TDATA = 50'b10101010000101111110101111011000111111101110010100;
        12'd2610: TDATA = 50'b10101010000011111001010101011000111100011100111100;
        12'd2611: TDATA = 50'b10101010000001110011110111011000111001001011100110;
        12'd2612: TDATA = 50'b10101001111111101110100111011000110101111010100111;
        12'd2613: TDATA = 50'b10101001111101101001011001011000110010101001110010;
        12'd2614: TDATA = 50'b10101001111011100100010001011000101111011001001100;
        12'd2615: TDATA = 50'b10101001111001011111001011011000101100001000101111;
        12'd2616: TDATA = 50'b10101001110111011010001001011000101000111000011100;
        12'd2617: TDATA = 50'b10101001110101010101010001011000100101101000011101;
        12'd2618: TDATA = 50'b10101001110011010000011011011000100010011000100111;
        12'd2619: TDATA = 50'b10101001110001001011101011011000011111001001000000;
        12'd2620: TDATA = 50'b10101001101111000110111011011000011011111001011101;
        12'd2621: TDATA = 50'b10101001101101000010010011011000011000101010001110;
        12'd2622: TDATA = 50'b10101001101010111101110011011000010101011011001101;
        12'd2623: TDATA = 50'b10101001101000111001010101011000010010001100010110;
        12'd2624: TDATA = 50'b10101001100110110100111101011000001110111101101110;
        12'd2625: TDATA = 50'b10101001100100110000100111011000001011101111001111;
        12'd2626: TDATA = 50'b10101001100010101100010011011000001000100000110101;
        12'd2627: TDATA = 50'b10101001100000101000001101011000000101010010111000;
        12'd2628: TDATA = 50'b10101001011110100100001001011000000010000101000100;
        12'd2629: TDATA = 50'b10101001011100100000000111010111111110110111010101;
        12'd2630: TDATA = 50'b10101001011010011100001001010111111011101001110101;
        12'd2631: TDATA = 50'b10101001011000011000011001010111111000011100101100;
        12'd2632: TDATA = 50'b10101001010110010100100001010111110101001111011111;
        12'd2633: TDATA = 50'b10101001010100010000110011010111110010000010100101;
        12'd2634: TDATA = 50'b10101001010010001101001011010111101110110101111001;
        12'd2635: TDATA = 50'b10101001010000001001100111010111101011101001010111;
        12'd2636: TDATA = 50'b10101001001110000110001011010111101000011101001000;
        12'd2637: TDATA = 50'b10101001001100000010110001010111100101010001000011;
        12'd2638: TDATA = 50'b10101001001001111111011001010111100010000101000010;
        12'd2639: TDATA = 50'b10101001000111111100001001010111011110111001010100;
        12'd2640: TDATA = 50'b10101001000101111000111111010111011011101101110101;
        12'd2641: TDATA = 50'b10101001000011110101110101010111011000100010011010;
        12'd2642: TDATA = 50'b10101001000001110010110011010111010101010111010011;
        12'd2643: TDATA = 50'b10101000111111101111111001010111010010001100011001;
        12'd2644: TDATA = 50'b10101000111101101100111011010111001111000001100000;
        12'd2645: TDATA = 50'b10101000111011101010001001010111001011110110111111;
        12'd2646: TDATA = 50'b10101000111001100111011001010111001000101100100111;
        12'd2647: TDATA = 50'b10101000110111100100101011010111000101100010010011;
        12'd2648: TDATA = 50'b10101000110101100010000111010111000010011000011000;
        12'd2649: TDATA = 50'b10101000110011011111100101010110111111001110100001;
        12'd2650: TDATA = 50'b10101000110001011101000111010110111100000100111000;
        12'd2651: TDATA = 50'b10101000101111011010110011010110111000111011100010;
        12'd2652: TDATA = 50'b10101000101101011000011101010110110101110010001100;
        12'd2653: TDATA = 50'b10101000101011010110010001010110110010101001001110;
        12'd2654: TDATA = 50'b10101000101001010100001001010110101111100000011001;
        12'd2655: TDATA = 50'b10101000100111010010000001010110101100010111101001;
        12'd2656: TDATA = 50'b10101000100101010000000011010110101001001111001100;
        12'd2657: TDATA = 50'b10101000100011001110000111010110100110000110111000;
        12'd2658: TDATA = 50'b10101000100001001100010001010110100010111110110010;
        12'd2659: TDATA = 50'b10101000011111001010100001010110011111110110111010;
        12'd2660: TDATA = 50'b10101000011101001000110001010110011100101111001000;
        12'd2661: TDATA = 50'b10101000011011000111001001010110011001100111100111;
        12'd2662: TDATA = 50'b10101000011001000101100011010110010110100000001100;
        12'd2663: TDATA = 50'b10101000010111000100000101010110010011011001000011;
        12'd2664: TDATA = 50'b10101000010101000010101101010110010000010010001000;
        12'd2665: TDATA = 50'b10101000010011000001010101010110001101001011010010;
        12'd2666: TDATA = 50'b10101000010000111111111111010110001010000100100110;
        12'd2667: TDATA = 50'b10101000001110111110111001010110000110111110010101;
        12'd2668: TDATA = 50'b10101000001100111101101011010110000011110111111011;
        12'd2669: TDATA = 50'b10101000001010111100100111010110000000110001111000;
        12'd2670: TDATA = 50'b10101000001000111011100111010101111101101011111111;
        12'd2671: TDATA = 50'b10101000000110111010110011010101111010100110011100;
        12'd2672: TDATA = 50'b10101000000100111001111001010101110111100000110110;
        12'd2673: TDATA = 50'b10101000000010111001001011010101110100011011100110;
        12'd2674: TDATA = 50'b10101000000000111000100001010101110001010110100000;
        12'd2675: TDATA = 50'b10100111111110110111111001010101101110010001100011;
        12'd2676: TDATA = 50'b10100111111100110111010011010101101011001100101111;
        12'd2677: TDATA = 50'b10100111111010110110110111010101101000001000001110;
        12'd2678: TDATA = 50'b10100111111000110110011001010101100101000011101101;
        12'd2679: TDATA = 50'b10100111110110110110000011010101100001111111011110;
        12'd2680: TDATA = 50'b10100111110100110101110011010101011110111011011110;
        12'd2681: TDATA = 50'b10100111110010110101100011010101011011110111100010;
        12'd2682: TDATA = 50'b10100111110000110101100001010101011000110100000001;
        12'd2683: TDATA = 50'b10100111101110110101100001010101010101110000100101;
        12'd2684: TDATA = 50'b10100111101100110101011111010101010010101101001110;
        12'd2685: TDATA = 50'b10100111101010110101100101010101001111101010000101;
        12'd2686: TDATA = 50'b10100111101000110101110011010101001100100111001110;
        12'd2687: TDATA = 50'b10100111100110110110000001010101001001100100011011;
        12'd2688: TDATA = 50'b10100111100100110110010001010101000110100001110010;
        12'd2689: TDATA = 50'b10100111100010110110101111010101000011011111100000;
        12'd2690: TDATA = 50'b10100111100000110111001011010101000000011101010010;
        12'd2691: TDATA = 50'b10100111011110110111101011010100111101011011001110;
        12'd2692: TDATA = 50'b10100111011100111000010001010100111010011001010111;
        12'd2693: TDATA = 50'b10100111011010111001000001010100110111010111110011;
        12'd2694: TDATA = 50'b10100111011000111001101001010100110100010110001010;
        12'd2695: TDATA = 50'b10100111010110111010100001010100110001010100111100;
        12'd2696: TDATA = 50'b10100111010100111011011001010100101110010011110011;
        12'd2697: TDATA = 50'b10100111010010111100010001010100101011010010101111;
        12'd2698: TDATA = 50'b10100111010000111101011001010100101000010010000110;
        12'd2699: TDATA = 50'b10100111001110111110011001010100100101010001011001;
        12'd2700: TDATA = 50'b10100111001100111111100111010100100010010001000010;
        12'd2701: TDATA = 50'b10100111001011000000110111010100011111010000110100;
        12'd2702: TDATA = 50'b10100111001001000010000111010100011100010000101011;
        12'd2703: TDATA = 50'b10100111000111000011100011010100011001010000111001;
        12'd2704: TDATA = 50'b10100111000101000100111011010100010110010001000110;
        12'd2705: TDATA = 50'b10100111000011000110011011010100010011010001100010;
        12'd2706: TDATA = 50'b10100111000001000111111111010100010000010010001011;
        12'd2707: TDATA = 50'b10100110111111001001101011010100001101010011000001;
        12'd2708: TDATA = 50'b10100110111101001011011011010100001010010100000101;
        12'd2709: TDATA = 50'b10100110111011001101001101010100000111010101001110;
        12'd2710: TDATA = 50'b10100110111001001111000111010100000100010110101000;
        12'd2711: TDATA = 50'b10100110110111010001000011010100000001011000001100;
        12'd2712: TDATA = 50'b10100110110101010011000011010011111110011001111001;
        12'd2713: TDATA = 50'b10100110110011010101000111010011111011011011101111;
        12'd2714: TDATA = 50'b10100110110001010111001001010011111000011101101001;
        12'd2715: TDATA = 50'b10100110101111011001011011010011110101011111111110;
        12'd2716: TDATA = 50'b10100110101101011011110001010011110010100010011100;
        12'd2717: TDATA = 50'b10100110101011011110001001010011101111100101000100;
        12'd2718: TDATA = 50'b10100110101001100000100001010011101100100111110000;
        12'd2719: TDATA = 50'b10100110100111100010111111010011101001101010101001;
        12'd2720: TDATA = 50'b10100110100101100101100011010011100110101101110000;
        12'd2721: TDATA = 50'b10100110100011101000001001010011100011110000111111;
        12'd2722: TDATA = 50'b10100110100001101010110111010011100000110100011101;
        12'd2723: TDATA = 50'b10100110011111101101100111010011011101111000000011;
        12'd2724: TDATA = 50'b10100110011101110000011101010011011010111011110110;
        12'd2725: TDATA = 50'b10100110011011110011010011010011010111111111101110;
        12'd2726: TDATA = 50'b10100110011001110110010101010011010101000011111101;
        12'd2727: TDATA = 50'b10100110010111111001011001010011010010001000010100;
        12'd2728: TDATA = 50'b10100110010101111100011111010011001111001100110000;
        12'd2729: TDATA = 50'b10100110010011111111101001010011001100010001011001;
        12'd2730: TDATA = 50'b10100110010010000010111011010011001001010110010000;
        12'd2731: TDATA = 50'b10100110010000000110001111010011000110011011001111;
        12'd2732: TDATA = 50'b10100110001110001001101001010011000011100000011100;
        12'd2733: TDATA = 50'b10100110001100001100111111010011000000100101101001;
        12'd2734: TDATA = 50'b10100110001010010000100011010010111101101011001100;
        12'd2735: TDATA = 50'b10100110001000010100001011010010111010110000111100;
        12'd2736: TDATA = 50'b10100110000110010111110101010010110111110110110001;
        12'd2737: TDATA = 50'b10100110000100011011100001010010110100111100101111;
        12'd2738: TDATA = 50'b10100110000010011111011001010010110010000011000010;
        12'd2739: TDATA = 50'b10100110000000100011001011010010101111001001010010;
        12'd2740: TDATA = 50'b10100101111110100111001011010010101100001111111100;
        12'd2741: TDATA = 50'b10100101111100101011001001010010101001010110100110;
        12'd2742: TDATA = 50'b10100101111010101111010001010010100110011101100001;
        12'd2743: TDATA = 50'b10100101111000110011010101010010100011100100011101;
        12'd2744: TDATA = 50'b10100101110110110111011111010010100000101011100110;
        12'd2745: TDATA = 50'b10100101110100111011110001010010011101110011000000;
        12'd2746: TDATA = 50'b10100101110011000000001011010010011010111010101000;
        12'd2747: TDATA = 50'b10100101110001000100100001010010011000000010010000;
        12'd2748: TDATA = 50'b10100101101111001000111111010010010101001010001001;
        12'd2749: TDATA = 50'b10100101101101001101100101010010010010010010001111;
        12'd2750: TDATA = 50'b10100101101011010010001001010010001111011010011010;
        12'd2751: TDATA = 50'b10100101101001010110110101010010001100100010110010;
        12'd2752: TDATA = 50'b10100101100111011011011111010010001001101011001110;
        12'd2753: TDATA = 50'b10100101100101100000011001010010000110110100000101;
        12'd2754: TDATA = 50'b10100101100011100101001011010010000011111100110011;
        12'd2755: TDATA = 50'b10100101100001101010000111010010000001000101110111;
        12'd2756: TDATA = 50'b10100101011111101111000111010001111110001111000011;
        12'd2757: TDATA = 50'b10100101011101110100010011010001111011011000100110;
        12'd2758: TDATA = 50'b10100101011011111001011001010001111000100010000100;
        12'd2759: TDATA = 50'b10100101011001111110101001010001110101101011110011;
        12'd2760: TDATA = 50'b10100101011000000011110111010001110010110101100111;
        12'd2761: TDATA = 50'b10100101010110001001001101010001101111111111101000;
        12'd2762: TDATA = 50'b10100101010100001110101011010001101101001001111010;
        12'd2763: TDATA = 50'b10100101010010010100001001010001101010010100010001;
        12'd2764: TDATA = 50'b10100101010000011001101001010001100111011110110001;
        12'd2765: TDATA = 50'b10100101001110011111010001010001100100101001011101;
        12'd2766: TDATA = 50'b10100101001100100100111011010001100001110100010010;
        12'd2767: TDATA = 50'b10100101001010101010101011010001011110111111010100;
        12'd2768: TDATA = 50'b10100101001000110000011011010001011100001010011010;
        12'd2769: TDATA = 50'b10100101000110110110010111010001011001010101110110;
        12'd2770: TDATA = 50'b10100101000100111100001111010001010110100001010010;
        12'd2771: TDATA = 50'b10100101000011000010010001010001010011101101000000;
        12'd2772: TDATA = 50'b10100101000001001000011001010001010000111000111010;
        12'd2773: TDATA = 50'b10100100111111001110100001010001001110000100111001;
        12'd2774: TDATA = 50'b10100100111101010100101101010001001011010001000000;
        12'd2775: TDATA = 50'b10100100111011011010111011010001001000011101010000;
        12'd2776: TDATA = 50'b10100100111001100001010001010001000101101001110001;
        12'd2777: TDATA = 50'b10100100110111100111101111010001000010110110011111;
        12'd2778: TDATA = 50'b10100100110101101110001011010001000000000011010010;
        12'd2779: TDATA = 50'b10100100110011110100101111010000111101010000010001;
        12'd2780: TDATA = 50'b10100100110001111011010101010000111010011101011001;
        12'd2781: TDATA = 50'b10100100110000000010000001010000110111101010101110;
        12'd2782: TDATA = 50'b10100100101110001000101101010000110100111000000110;
        12'd2783: TDATA = 50'b10100100101100001111100001010000110010000101110001;
        12'd2784: TDATA = 50'b10100100101010010110010111010000101111010011011111;
        12'd2785: TDATA = 50'b10100100101000011101010001010000101100100001011010;
        12'd2786: TDATA = 50'b10100100100110100100001111010000101001101111011110;
        12'd2787: TDATA = 50'b10100100100100101011010111010000100110111101110011;
        12'd2788: TDATA = 50'b10100100100010110010100001010000100100001100010001;
        12'd2789: TDATA = 50'b10100100100000111001100101010000100001011010101010;
        12'd2790: TDATA = 50'b10100100011111000000110111010000011110101001011100;
        12'd2791: TDATA = 50'b10100100011101001000001011010000011011111000010011;
        12'd2792: TDATA = 50'b10100100011011001111100011010000011001000111010111;
        12'd2793: TDATA = 50'b10100100011001010111000011010000010110010110101000;
        12'd2794: TDATA = 50'b10100100010111011110100101010000010011100110000001;
        12'd2795: TDATA = 50'b10100100010101100110000111010000010000110101011110;
        12'd2796: TDATA = 50'b10100100010011101101110001010000001110000101001101;
        12'd2797: TDATA = 50'b10100100010001110101011001010000001011010100111011;
        12'd2798: TDATA = 50'b10100100001111111101001011010000001000100100111010;
        12'd2799: TDATA = 50'b10100100001110000101000001010000000101110101000110;
        12'd2800: TDATA = 50'b10100100001100001100111011010000000011000101011011;
        12'd2801: TDATA = 50'b10100100001010010100111011010000000000010101111100;
        12'd2802: TDATA = 50'b10100100001000011100111011001111111101100110100001;
        12'd2803: TDATA = 50'b10100100000110100100111111001111111010110111001111;
        12'd2804: TDATA = 50'b10100100000100101101000111001111111000001000001001;
        12'd2805: TDATA = 50'b10100100000010110101010111001111110101011001010000;
        12'd2806: TDATA = 50'b10100100000000111101101011001111110010101010100100;
        12'd2807: TDATA = 50'b10100011111111000110000001001111101111111011111100;
        12'd2808: TDATA = 50'b10100011111101001110011001001111101101001101011101;
        12'd2809: TDATA = 50'b10100011111011010110110111001111101010011111001010;
        12'd2810: TDATA = 50'b10100011111001011111011011001111100111110001000011;
        12'd2811: TDATA = 50'b10100011110111101000000001001111100101000011000101;
        12'd2812: TDATA = 50'b10100011110101110000101001001111100010010101001011;
        12'd2813: TDATA = 50'b10100011110011111001011001001111011111100111100010;
        12'd2814: TDATA = 50'b10100011110010000010001111001111011100111010000110;
        12'd2815: TDATA = 50'b10100011110000001011000001001111011010001100101001;
        12'd2816: TDATA = 50'b10100011101110010011111011001111010111011111011001;
        12'd2817: TDATA = 50'b10100011101100011100111101001111010100110010011011;
        12'd2818: TDATA = 50'b10100011101010100110000001001111010010000101100100;
        12'd2819: TDATA = 50'b10100011101000101111000111001111001111011000110001;
        12'd2820: TDATA = 50'b10100011100110111000010001001111001100101100001011;
        12'd2821: TDATA = 50'b10100011100101000001011111001111001001111111101101;
        12'd2822: TDATA = 50'b10100011100011001010110011001111000111010011011100;
        12'd2823: TDATA = 50'b10100011100001010100001011001111000100100111010011;
        12'd2824: TDATA = 50'b10100011011111011101100101001111000001111011010010;
        12'd2825: TDATA = 50'b10100011011101100111000101001110111111001111011110;
        12'd2826: TDATA = 50'b10100011011011110000100101001110111100100011101110;
        12'd2827: TDATA = 50'b10100011011001111010010001001110111001111000010011;
        12'd2828: TDATA = 50'b10100011011000000011111001001110110111001100110111;
        12'd2829: TDATA = 50'b10100011010110001101101001001110110100100001101001;
        12'd2830: TDATA = 50'b10100011010100010111011011001110110001110110100010;
        12'd2831: TDATA = 50'b10100011010010100001010011001110101111001011101000;
        12'd2832: TDATA = 50'b10100011010000101011001011001110101100100000110010;
        12'd2833: TDATA = 50'b10100011001110110101001111001110101001110110010000;
        12'd2834: TDATA = 50'b10100011001100111111001111001110100111001011101111;
        12'd2835: TDATA = 50'b10100011001011001001010111001110100100100001011010;
        12'd2836: TDATA = 50'b10100011001001010011100001001110100001110111001101;
        12'd2837: TDATA = 50'b10100011000111011101110001001110011111001101001101;
        12'd2838: TDATA = 50'b10100011000101101000000111001110011100100011011001;
        12'd2839: TDATA = 50'b10100011000011110010011101001110011001111001101001;
        12'd2840: TDATA = 50'b10100011000001111100111001001110010111010000000110;
        12'd2841: TDATA = 50'b10100011000000000111010111001110010100100110101010;
        12'd2842: TDATA = 50'b10100010111110010001111101001110010001111101011011;
        12'd2843: TDATA = 50'b10100010111100011100100001001110001111010100010000;
        12'd2844: TDATA = 50'b10100010111010100111001101001110001100101011010010;
        12'd2845: TDATA = 50'b10100010111000110001110111001110001010000010010111;
        12'd2846: TDATA = 50'b10100010110110111100110001001110000111011001110101;
        12'd2847: TDATA = 50'b10100010110101000111100011001110000100110001001011;
        12'd2848: TDATA = 50'b10100010110011010010011111001110000010001000110101;
        12'd2849: TDATA = 50'b10100010110001011101011101001101111111100000100011;
        12'd2850: TDATA = 50'b10100010101111101000011111001101111100111000011110;
        12'd2851: TDATA = 50'b10100010101101110011101011001101111010010000101001;
        12'd2852: TDATA = 50'b10100010101011111110110001001101110111101000110000;
        12'd2853: TDATA = 50'b10100010101010001010000011001101110101000001001011;
        12'd2854: TDATA = 50'b10100010101000010101011001001101110010011001101111;
        12'd2855: TDATA = 50'b10100010100110100000101011001101101111110010010010;
        12'd2856: TDATA = 50'b10100010100100101100001001001101101101001011001010;
        12'd2857: TDATA = 50'b10100010100010110111100001001101101010100011111101;
        12'd2858: TDATA = 50'b10100010100001000011000001001101100111111101000000;
        12'd2859: TDATA = 50'b10100010011111001110101001001101100101010110010000;
        12'd2860: TDATA = 50'b10100010011101011010010011001101100010101111101000;
        12'd2861: TDATA = 50'b10100010011011100110000011001101100000001001001101;
        12'd2862: TDATA = 50'b10100010011001110001110011001101011101100010110101;
        12'd2863: TDATA = 50'b10100010010111111101101001001101011010111100101001;
        12'd2864: TDATA = 50'b10100010010110001001100001001101011000010110100110;
        12'd2865: TDATA = 50'b10100010010100010101100001001101010101110000101111;
        12'd2866: TDATA = 50'b10100010010010100001011111001101010011001010111011;
        12'd2867: TDATA = 50'b10100010010000101101100101001101010000100101010100;
        12'd2868: TDATA = 50'b10100010001110111001101111001101001101111111111001;
        12'd2869: TDATA = 50'b10100010001101000101111011001101001011011010100001;
        12'd2870: TDATA = 50'b10100010001011010010001111001101001000110101011010;
        12'd2871: TDATA = 50'b10100010001001011110100011001101000110010000010111;
        12'd2872: TDATA = 50'b10100010000111101010111001001101000011101011011100;
        12'd2873: TDATA = 50'b10100010000101110111010111001101000001000110101101;
        12'd2874: TDATA = 50'b10100010000100000011110111001100111110100010000110;
        12'd2875: TDATA = 50'b10100010000010010000011101001100111011111101101011;
        12'd2876: TDATA = 50'b10100010000000011101000011001100111001011001010100;
        12'd2877: TDATA = 50'b10100001111110101001110001001100110110110101001101;
        12'd2878: TDATA = 50'b10100001111100110110100001001100110100010001001010;
        12'd2879: TDATA = 50'b10100001111011000011010011001100110001101101001111;
        12'd2880: TDATA = 50'b10100001111001010000000111001100101111001001011100;
        12'd2881: TDATA = 50'b10100001110111011101000011001100101100100101110101;
        12'd2882: TDATA = 50'b10100001110101101010000111001100101010000010011111;
        12'd2883: TDATA = 50'b10100001110011110111000101001100100111011111000011;
        12'd2884: TDATA = 50'b10100001110010000100001111001100100100111011111100;
        12'd2885: TDATA = 50'b10100001110000010001011001001100100010011000111001;
        12'd2886: TDATA = 50'b10100001101110011110101001001100011111110110000010;
        12'd2887: TDATA = 50'b10100001101100101011111001001100011101010011001110;
        12'd2888: TDATA = 50'b10100001101010111001001111001100011010110000100111;
        12'd2889: TDATA = 50'b10100001101001000110101011001100011000001110001100;
        12'd2890: TDATA = 50'b10100001100111010100000111001100010101101011110100;
        12'd2891: TDATA = 50'b10100001100101100001100011001100010011001001100000;
        12'd2892: TDATA = 50'b10100001100011101111001011001100010000100111100001;
        12'd2893: TDATA = 50'b10100001100001111100110011001100001110000101100101;
        12'd2894: TDATA = 50'b10100001100000001010100011001100001011100011111001;
        12'd2895: TDATA = 50'b10100001011110011000010001001100001001000010001101;
        12'd2896: TDATA = 50'b10100001011100100110000011001100000110100000101000;
        12'd2897: TDATA = 50'b10100001011010110011111101001100000011111111010100;
        12'd2898: TDATA = 50'b10100001011001000001111101001100000001011110001100;
        12'd2899: TDATA = 50'b10100001010111001111111001001011111110111101000100;
        12'd2900: TDATA = 50'b10100001010101011101111101001011111100011100000111;
        12'd2901: TDATA = 50'b10100001010011101100001001001011111001111011011010;
        12'd2902: TDATA = 50'b10100001010001111010010001001011110111011010101101;
        12'd2903: TDATA = 50'b10100001010000001000100001001011110100111010001100;
        12'd2904: TDATA = 50'b10100001001110010110110011001011110010011001110011;
        12'd2905: TDATA = 50'b10100001001100100101001011001011101111111001100101;
        12'd2906: TDATA = 50'b10100001001010110011100011001011101101011001011011;
        12'd2907: TDATA = 50'b10100001001001000010000001001011101010111001011101;
        12'd2908: TDATA = 50'b10100001000111010000100001001011101000011001100111;
        12'd2909: TDATA = 50'b10100001000101011111001001001011100101111001111101;
        12'd2910: TDATA = 50'b10100001000011101101101111001011100011011010010110;
        12'd2911: TDATA = 50'b10100001000001111100011101001011100000111010111100;
        12'd2912: TDATA = 50'b10100001000000001011001101001011011110011011101001;
        12'd2913: TDATA = 50'b10100000111110011010000011001011011011111100100010;
        12'd2914: TDATA = 50'b10100000111100101000111001001011011001011101011110;
        12'd2915: TDATA = 50'b10100000111010110111110101001011010110111110100110;
        12'd2916: TDATA = 50'b10100000111001000110110011001011010100011111110111;
        12'd2917: TDATA = 50'b10100000110111010101111001001011010010000001010011;
        12'd2918: TDATA = 50'b10100000110101100101000001001011001111100010110110;
        12'd2919: TDATA = 50'b10100000110011110100001001001011001101000100011101;
        12'd2920: TDATA = 50'b10100000110010000011010111001011001010100110010000;
        12'd2921: TDATA = 50'b10100000110000010010101011001011001000001000001111;
        12'd2922: TDATA = 50'b10100000101110100001111111001011000101101010010010;
        12'd2923: TDATA = 50'b10100000101100110001011011001011000011001100100100;
        12'd2924: TDATA = 50'b10100000101011000000110011001011000000101110110001;
        12'd2925: TDATA = 50'b10100000101001010000011001001010111110010001011000;
        12'd2926: TDATA = 50'b10100000100111011111111011001010111011110011111101;
        12'd2927: TDATA = 50'b10100000100101101111100001001010111001010110101001;
        12'd2928: TDATA = 50'b10100000100011111111010001001010110110111001100110;
        12'd2929: TDATA = 50'b10100000100010001110111101001010110100011100100010;
        12'd2930: TDATA = 50'b10100000100000011110110001001010110001111111101111;
        12'd2931: TDATA = 50'b10100000011110101110101001001010101111100011000010;
        12'd2932: TDATA = 50'b10100000011100111110100001001010101101000110011001;
        12'd2933: TDATA = 50'b10100000011011001110011111001010101010101001111100;
        12'd2934: TDATA = 50'b10100000011001011110100011001010101000001101101011;
        12'd2935: TDATA = 50'b10100000010111101110100111001010100101110001011101;
        12'd2936: TDATA = 50'b10100000010101111110101111001010100011010101010111;
        12'd2937: TDATA = 50'b10100000010100001110111111001010100000111001100001;
        12'd2938: TDATA = 50'b10100000010010011111001111001010011110011101101110;
        12'd2939: TDATA = 50'b10100000010000101111100001001010011100000010000010;
        12'd2940: TDATA = 50'b10100000001110111111111011001010011001100110100011;
        12'd2941: TDATA = 50'b10100000001101010000010011001010010111001011000110;
        12'd2942: TDATA = 50'b10100000001011100000110011001010010100101111110110;
        12'd2943: TDATA = 50'b10100000001001110001010111001010010010010100110001;
        12'd2944: TDATA = 50'b10100000001000000001111111001010001111111001110100;
        12'd2945: TDATA = 50'b10100000000110010010100111001010001101011110111010;
        12'd2946: TDATA = 50'b10100000000100100011010011001010001011000100001000;
        12'd2947: TDATA = 50'b10100000000010110100001001001010001000101001101010;
        12'd2948: TDATA = 50'b10100000000001000100110111001010000110001111000010;
        12'd2949: TDATA = 50'b10011111111111010101110101001010000011110100110011;
        12'd2950: TDATA = 50'b10011111111101100110110001001010000001011010100111;
        12'd2951: TDATA = 50'b10011111111011110111101111001001111111000000011110;
        12'd2952: TDATA = 50'b10011111111010001000110001001001111100100110100010;
        12'd2953: TDATA = 50'b10011111111000011001110111001001111010001100101100;
        12'd2954: TDATA = 50'b10011111110110101011000111001001110111110011000111;
        12'd2955: TDATA = 50'b10011111110100111100010011001001110101011001100000;
        12'd2956: TDATA = 50'b10011111110011001101100001001001110011000000000001;
        12'd2957: TDATA = 50'b10011111110001011110110111001001110000100110101110;
        12'd2958: TDATA = 50'b10011111101111110000001111001001101110001101100010;
        12'd2959: TDATA = 50'b10011111101110000001101111001001101011110100100110;
        12'd2960: TDATA = 50'b10011111101100010011010001001001101001011011101101;
        12'd2961: TDATA = 50'b10011111101010100100110001001001100111000010111000;
        12'd2962: TDATA = 50'b10011111101000110110011001001001100100101010001110;
        12'd2963: TDATA = 50'b10011111100111001000000011001001100010010001101100;
        12'd2964: TDATA = 50'b10011111100101011001110011001001011111111001010101;
        12'd2965: TDATA = 50'b10011111100011101011100011001001011101100001000001;
        12'd2966: TDATA = 50'b10011111100001111101011011001001011011001000111110;
        12'd2967: TDATA = 50'b10011111100000001111010101001001011000110000111101;
        12'd2968: TDATA = 50'b10011111011110100001010001001001010110011001000100;
        12'd2969: TDATA = 50'b10011111011100110011001111001001010100000001010010;
        12'd2970: TDATA = 50'b10011111011011000101010001001001010001101001101000;
        12'd2971: TDATA = 50'b10011111011001010111011001001001001111010010001001;
        12'd2972: TDATA = 50'b10011111010111101001100101001001001100111010110010;
        12'd2973: TDATA = 50'b10011111010101111011110011001001001010100011100010;
        12'd2974: TDATA = 50'b10011111010100001110000111001001001000001100011110;
        12'd2975: TDATA = 50'b10011111010010100000011011001001000101110101011100;
        12'd2976: TDATA = 50'b10011111010000110010110101001001000011011110100111;
        12'd2977: TDATA = 50'b10011111001111000101001111001001000001000111110100;
        12'd2978: TDATA = 50'b10011111001101010111110001001000111110110001010001;
        12'd2979: TDATA = 50'b10011111001011101010010101001000111100011010110010;
        12'd2980: TDATA = 50'b10011111001001111100111011001000111010000100011010;
        12'd2981: TDATA = 50'b10011111001000001111101001001000110111101110010001;
        12'd2982: TDATA = 50'b10011111000110100010011001001000110101011000001100;
        12'd2983: TDATA = 50'b10011111000100110101000101001000110011000010000101;
        12'd2984: TDATA = 50'b10011111000011000111111001001000110000101100001111;
        12'd2985: TDATA = 50'b10011111000001011010110001001000101110010110011111;
        12'd2986: TDATA = 50'b10011110111111101101101111001000101100000000111011;
        12'd2987: TDATA = 50'b10011110111110000000110011001000101001101011100011;
        12'd2988: TDATA = 50'b10011110111100010011110001001000100111010110000101;
        12'd2989: TDATA = 50'b10011110111010100110111011001000100101000000111011;
        12'd2990: TDATA = 50'b10011110111000111010001001001000100010101011111001;
        12'd2991: TDATA = 50'b10011110110111001101010011001000100000010110110101;
        12'd2992: TDATA = 50'b10011110110101100000100011001000011110000001111101;
        12'd2993: TDATA = 50'b10011110110011110011111001001000011011101101010000;
        12'd2994: TDATA = 50'b10011110110010000111010001001000011001011000101011;
        12'd2995: TDATA = 50'b10011110110000011010101011001000010111000100001001;
        12'd2996: TDATA = 50'b10011110101110101110001101001000010100101111110110;
        12'd2997: TDATA = 50'b10011110101101000001101111001000010010011011100110;
        12'd2998: TDATA = 50'b10011110101011010101010111001000010000000111100010;
        12'd2999: TDATA = 50'b10011110101001101001000001001000001101110011100101;
        12'd3000: TDATA = 50'b10011110100111111100101001001000001011011111100111;
        12'd3001: TDATA = 50'b10011110100110010000010111001000001001001011110100;
        12'd3002: TDATA = 50'b10011110100100100100010001001000000110111000010101;
        12'd3003: TDATA = 50'b10011110100010111000000011001000000100100100101101;
        12'd3004: TDATA = 50'b10011110100001001011111111001000000010010001011000;
        12'd3005: TDATA = 50'b10011110011111011111111111000111111111111110001011;
        12'd3006: TDATA = 50'b10011110011101110011111111000111111101101011000000;
        12'd3007: TDATA = 50'b10011110011100001000001011000111111011011000001010;
        12'd3008: TDATA = 50'b10011110011010011100001111000111111001000101001010;
        12'd3009: TDATA = 50'b10011110011000110000100001000111110110110010100001;
        12'd3010: TDATA = 50'b10011110010111000100101001000111110100011111101111;
        12'd3011: TDATA = 50'b10011110010101011000111111000111110010001101010001;
        12'd3012: TDATA = 50'b10011110010011101101010011000111101111111010110110;
        12'd3013: TDATA = 50'b10011110010010000001101011000111101101101000100010;
        12'd3014: TDATA = 50'b10011110010000010110001101000111101011010110011110;
        12'd3015: TDATA = 50'b10011110001110101010110001000111101001000100100001;
        12'd3016: TDATA = 50'b10011110001100111111010001000111100110110010100010;
        12'd3017: TDATA = 50'b10011110001011010011111001000111100100100000101111;
        12'd3018: TDATA = 50'b10011110001001101000100011000111100010001111000011;
        12'd3019: TDATA = 50'b10011110000111111101010011000111011111111101100011;
        12'd3020: TDATA = 50'b10011110000110010010000011000111011101101100000101;
        12'd3021: TDATA = 50'b10011110000100100110110011000111011011011010101011;
        12'd3022: TDATA = 50'b10011110000010111011110001000111011001001001101000;
        12'd3023: TDATA = 50'b10011110000001010000101011000111010110111000011111;
        12'd3024: TDATA = 50'b10011101111111100101101101000111010100100111100111;
        12'd3025: TDATA = 50'b10011101111101111010110001000111010010010110110101;
        12'd3026: TDATA = 50'b10011101111100001111110111000111010000000110000110;
        12'd3027: TDATA = 50'b10011101111010100100111111000111001101110101011110;
        12'd3028: TDATA = 50'b10011101111000111010001001000111001011100100111110;
        12'd3029: TDATA = 50'b10011101110111001111011011000111001001010100101001;
        12'd3030: TDATA = 50'b10011101110101100100101111000111000111000100011011;
        12'd3031: TDATA = 50'b10011101110011111010000011000111000100110100001111;
        12'd3032: TDATA = 50'b10011101110010001111011111000111000010100100010011;
        12'd3033: TDATA = 50'b10011101110000100100111101000111000000010100011010;
        12'd3034: TDATA = 50'b10011101101110111010011111000110111110000100101101;
        12'd3035: TDATA = 50'b10011101101101010000000011000110111011110101000010;
        12'd3036: TDATA = 50'b10011101101011100101101011000110111001100101100010;
        12'd3037: TDATA = 50'b10011101101001111011010101000110110111010110000110;
        12'd3038: TDATA = 50'b10011101101000010001000111000110110101000110111000;
        12'd3039: TDATA = 50'b10011101100110100110111001000110110010110111101110;
        12'd3040: TDATA = 50'b10011101100100111100110001000110110000101000101111;
        12'd3041: TDATA = 50'b10011101100011010010101001000110101110011001110010;
        12'd3042: TDATA = 50'b10011101100001101000100011000110101100001010111101;
        12'd3043: TDATA = 50'b10011101011111111110100001000110101001111100001111;
        12'd3044: TDATA = 50'b10011101011110010100101001000110100111101101110000;
        12'd3045: TDATA = 50'b10011101011100101010101001000110100101011111001011;
        12'd3046: TDATA = 50'b10011101011011000000110111000110100011010000111010;
        12'd3047: TDATA = 50'b10011101011001010111000001000110100001000010101000;
        12'd3048: TDATA = 50'b10011101010111101101010001000110011110110100100001;
        12'd3049: TDATA = 50'b10011101010110000011100111000110011100100110100101;
        12'd3050: TDATA = 50'b10011101010100011001111001000110011010011000101000;
        12'd3051: TDATA = 50'b10011101010010110000010011000110011000001010110110;
        12'd3052: TDATA = 50'b10011101010001000110110101000110010101111101010011;
        12'd3053: TDATA = 50'b10011101001111011101010001000110010011101111101011;
        12'd3054: TDATA = 50'b10011101001101110011110011000110010001100010001110;
        12'd3055: TDATA = 50'b10011101001100001010011011000110001111010100111100;
        12'd3056: TDATA = 50'b10011101001010100001001001000110001101000111110101;
        12'd3057: TDATA = 50'b10011101001000110111111001000110001010111010110101;
        12'd3058: TDATA = 50'b10011101000111001110100111000110001000101101110100;
        12'd3059: TDATA = 50'b10011101000101100101100001000110000110100001000110;
        12'd3060: TDATA = 50'b10011101000011111100010011000110000100010100001110;
        12'd3061: TDATA = 50'b10011101000010010011001111000110000010000111101010;
        12'd3062: TDATA = 50'b10011101000000101010001101000101111111111011001001;
        12'd3063: TDATA = 50'b10011100111111000001001111000101111101101110110011;
        12'd3064: TDATA = 50'b10011100111101011000011001000101111011100010100111;
        12'd3065: TDATA = 50'b10011100111011101111011111000101111001010110011011;
        12'd3066: TDATA = 50'b10011100111010000110100111000101110111001010010101;
        12'd3067: TDATA = 50'b10011100111000011101111001000101110100111110011111;
        12'd3068: TDATA = 50'b10011100110110110101001011000101110010110010101011;
        12'd3069: TDATA = 50'b10011100110101001100100001000101110000100110111110;
        12'd3070: TDATA = 50'b10011100110011100011111001000101101110011011011001;
        12'd3071: TDATA = 50'b10011100110001111011010011000101101100001111111010;
        12'd3072: TDATA = 50'b10011100110000010010110101000101101010000100100110;
        12'd3073: TDATA = 50'b10011100101110101010011001000101100111111001011001;
        12'd3074: TDATA = 50'b10011100101101000001111101000101100101101110001110;
        12'd3075: TDATA = 50'b10011100101011011001100111000101100011100011001111;
        12'd3076: TDATA = 50'b10011100101001110001010001000101100001011000010011;
        12'd3077: TDATA = 50'b10011100101000001001000001000101011111001101100001;
        12'd3078: TDATA = 50'b10011100100110100000110111000101011101000010111010;
        12'd3079: TDATA = 50'b10011100100100111000101001000101011010111000010011;
        12'd3080: TDATA = 50'b10011100100011010000100011000101011000101101110110;
        12'd3081: TDATA = 50'b10011100100001101000100001000101010110100011100100;
        12'd3082: TDATA = 50'b10011100100000000000100001000101010100011001010100;
        12'd3083: TDATA = 50'b10011100011110011000011111000101010010001111001000;
        12'd3084: TDATA = 50'b10011100011100110000100111000101010000000101001011;
        12'd3085: TDATA = 50'b10011100011011001000110011000101001101111011010100;
        12'd3086: TDATA = 50'b10011100011001100001000001000101001011110001100100;
        12'd3087: TDATA = 50'b10011100010111111001001111000101001001100111110111;
        12'd3088: TDATA = 50'b10011100010110010001100011000101000111011110010101;
        12'd3089: TDATA = 50'b10011100010100101001111001000101000101010100111010;
        12'd3090: TDATA = 50'b10011100010011000010010011000101000011001011100101;
        12'd3091: TDATA = 50'b10011100010001011010110011000101000001000010011011;
        12'd3092: TDATA = 50'b10011100001111110011010001000100111110111001010001;
        12'd3093: TDATA = 50'b10011100001110001011110011000100111100110000010000;
        12'd3094: TDATA = 50'b10011100001100100100011001000100111010100111010111;
        12'd3095: TDATA = 50'b10011100001010111101000011000100111000011110100101;
        12'd3096: TDATA = 50'b10011100001001010101110001000100110110010101111101;
        12'd3097: TDATA = 50'b10011100000111101110100001000100110100001101011000;
        12'd3098: TDATA = 50'b10011100000110000111010011000100110010000100111010;
        12'd3099: TDATA = 50'b10011100000100100000000111000100101111111100100011;
        12'd3100: TDATA = 50'b10011100000010111001000011000100101101110100010110;
        12'd3101: TDATA = 50'b10011100000001010010000011000100101011101100010100;
        12'd3102: TDATA = 50'b10011011111111101011000001000100101001100100010010;
        12'd3103: TDATA = 50'b10011011111110000100000011000100100111011100010101;
        12'd3104: TDATA = 50'b10011011111100011101001001000100100101010100100100;
        12'd3105: TDATA = 50'b10011011111010110110010011000100100011001100111001;
        12'd3106: TDATA = 50'b10011011111001001111100001000100100001000101010101;
        12'd3107: TDATA = 50'b10011011110111101000110001000100011110111101111000;
        12'd3108: TDATA = 50'b10011011110110000010000011000100011100110110100001;
        12'd3109: TDATA = 50'b10011011110100011011011001000100011010101111010010;
        12'd3110: TDATA = 50'b10011011110010110100110011000100011000101000001001;
        12'd3111: TDATA = 50'b10011011110001001110010001000100010110100001001010;
        12'd3112: TDATA = 50'b10011011101111100111101011000100010100011010000111;
        12'd3113: TDATA = 50'b10011011101110000001010011000100010010010011011010;
        12'd3114: TDATA = 50'b10011011101100011010110111000100010000001100101100;
        12'd3115: TDATA = 50'b10011011101010110100011111000100001110000110000100;
        12'd3116: TDATA = 50'b10011011101001001110001011000100001011111111100100;
        12'd3117: TDATA = 50'b10011011100111101000000001000100001001111001010110;
        12'd3118: TDATA = 50'b10011011100110000001101111000100000111110010111110;
        12'd3119: TDATA = 50'b10011011100100011011101001000100000101101100111010;
        12'd3120: TDATA = 50'b10011011100010110101100011000100000011100110111000;
        12'd3121: TDATA = 50'b10011011100001001111010111000100000001100000110001;
        12'd3122: TDATA = 50'b10011011011111101001010111000011111111011010111100;
        12'd3123: TDATA = 50'b10011011011110000011100011000011111101010101011010;
        12'd3124: TDATA = 50'b10011011011100011101100011000011111011001111101011;
        12'd3125: TDATA = 50'b10011011011010110111101001000011111001001010000110;
        12'd3126: TDATA = 50'b10011011011001010001111011000011110111000100110100;
        12'd3127: TDATA = 50'b10011011010111101100000001000011110100111111010101;
        12'd3128: TDATA = 50'b10011011010110000110011001000011110010111010010000;
        12'd3129: TDATA = 50'b10011011010100100000101011000011110000110101000110;
        12'd3130: TDATA = 50'b10011011010010111011000011000011101110110000000111;
        12'd3131: TDATA = 50'b10011011010001010101011111000011101100101011001110;
        12'd3132: TDATA = 50'b10011011001111110000000011000011101010100110100100;
        12'd3133: TDATA = 50'b10011011001110001010100001000011101000100001110101;
        12'd3134: TDATA = 50'b10011011001100100101000111000011100110011101010100;
        12'd3135: TDATA = 50'b10011011001010111111110001000011100100011000111010;
        12'd3136: TDATA = 50'b10011011001001011010011001000011100010010100011110;
        12'd3137: TDATA = 50'b10011011000111110101001001000011100000010000010010;
        12'd3138: TDATA = 50'b10011011000110001111111001000011011110001100000111;
        12'd3139: TDATA = 50'b10011011000100101010101111000011011100001000000111;
        12'd3140: TDATA = 50'b10011011000011000101100101000011011010000100001010;
        12'd3141: TDATA = 50'b10011011000001100000011011000011011000000000010000;
        12'd3142: TDATA = 50'b10011010111111111011011101000011010101111100101000;
        12'd3143: TDATA = 50'b10011010111110010110011011000011010011111000111111;
        12'd3144: TDATA = 50'b10011010111100110001100001000011010001110101100000;
        12'd3145: TDATA = 50'b10011010111011001100101001000011001111110010001000;
        12'd3146: TDATA = 50'b10011010111001100111110001000011001101101110110010;
        12'd3147: TDATA = 50'b10011010111000000010111111000011001011101011100111;
        12'd3148: TDATA = 50'b10011010110110011110001101000011001001101000011111;
        12'd3149: TDATA = 50'b10011010110100111001100011000011000111100101100101;
        12'd3150: TDATA = 50'b10011010110011010100110111000011000101100010101010;
        12'd3151: TDATA = 50'b10011010110001110000001111000011000011011111110101;
        12'd3152: TDATA = 50'b10011010110000001011101111000011000001011101001110;
        12'd3153: TDATA = 50'b10011010101110100111001111000010111111011010101011;
        12'd3154: TDATA = 50'b10011010101101000010101111000010111101011000001010;
        12'd3155: TDATA = 50'b10011010101011011110010101000010111011010101110011;
        12'd3156: TDATA = 50'b10011010101001111010000001000010111001010011100111;
        12'd3157: TDATA = 50'b10011010101000010101101001000010110111010001011010;
        12'd3158: TDATA = 50'b10011010100110110001011001000010110101001111010111;
        12'd3159: TDATA = 50'b10011010100101001101000101000010110011001101010010;
        12'd3160: TDATA = 50'b10011010100011101000111101000010110001001011100000;
        12'd3161: TDATA = 50'b10011010100010000100110101000010101111001001110001;
        12'd3162: TDATA = 50'b10011010100000100000101111000010101101001000001000;
        12'd3163: TDATA = 50'b10011010011110111100101011000010101011000110100010;
        12'd3164: TDATA = 50'b10011010011101011000101111000010101001000101001010;
        12'd3165: TDATA = 50'b10011010011011110100110011000010100111000011110100;
        12'd3166: TDATA = 50'b10011010011010010000111001000010100101000010100101;
        12'd3167: TDATA = 50'b10011010011000101101000011000010100011000001011101;
        12'd3168: TDATA = 50'b10011010010111001001010001000010100001000000011011;
        12'd3169: TDATA = 50'b10011010010101100101100001000010011110111111011111;
        12'd3170: TDATA = 50'b10011010010100000001110011000010011100111110101010;
        12'd3171: TDATA = 50'b10011010010010011110001001000010011010111101111100;
        12'd3172: TDATA = 50'b10011010010000111010100011000010011000111101010100;
        12'd3173: TDATA = 50'b10011010001111010110111111000010010110111100110010;
        12'd3174: TDATA = 50'b10011010001101110011011011000010010100111100010011;
        12'd3175: TDATA = 50'b10011010001100001111111111000010010010111100000011;
        12'd3176: TDATA = 50'b10011010001010101100100101000010010000111011110100;
        12'd3177: TDATA = 50'b10011010001001001001001101000010001110111011101101;
        12'd3178: TDATA = 50'b10011010000111100101110111000010001100111011101011;
        12'd3179: TDATA = 50'b10011010000110000010100011000010001010111011101101;
        12'd3180: TDATA = 50'b10011010000100011111011001000010001000111100000000;
        12'd3181: TDATA = 50'b10011010000010111100000111000010000110111100001010;
        12'd3182: TDATA = 50'b10011010000001011001000001000010000100111100100111;
        12'd3183: TDATA = 50'b10011001111111110101111111000010000010111101001001;
        12'd3184: TDATA = 50'b10011001111110010010111011000010000000111101101111;
        12'd3185: TDATA = 50'b10011001111100101111111011000001111110111110011010;
        12'd3186: TDATA = 50'b10011001111011001100111111000001111100111111001101;
        12'd3187: TDATA = 50'b10011001111001101010000001000001111011000000000001;
        12'd3188: TDATA = 50'b10011001111000000111010001000001111001000001001000;
        12'd3189: TDATA = 50'b10011001110110100100010111000001110111000010000110;
        12'd3190: TDATA = 50'b10011001110101000001101001000001110101000011010101;
        12'd3191: TDATA = 50'b10011001110011011110110111000001110011000100100011;
        12'd3192: TDATA = 50'b10011001110001111100001101000001110001000101111100;
        12'd3193: TDATA = 50'b10011001110000011001100101000001101111000111011011;
        12'd3194: TDATA = 50'b10011001101110110111000011000001101101001001000100;
        12'd3195: TDATA = 50'b10011001101101010100100001000001101011001010110000;
        12'd3196: TDATA = 50'b10011001101011110001111111000001101001001100011110;
        12'd3197: TDATA = 50'b10011001101010001111100011000001100111001110010110;
        12'd3198: TDATA = 50'b10011001101000101101001001000001100101010000010101;
        12'd3199: TDATA = 50'b10011001100111001010110001000001100011010010010111;
        12'd3200: TDATA = 50'b10011001100101101000100001000001100001010100100110;
        12'd3201: TDATA = 50'b10011001100100000110010001000001011111010110111000;
        12'd3202: TDATA = 50'b10011001100010100100000001000001011101011001001100;
        12'd3203: TDATA = 50'b10011001100001000001110111000001011011011011101011;
        12'd3204: TDATA = 50'b10011001011111011111101101000001011001011110001100;
        12'd3205: TDATA = 50'b10011001011101111101101011000001010111100000111011;
        12'd3206: TDATA = 50'b10011001011100011011100101000001010101100011100101;
        12'd3207: TDATA = 50'b10011001011010111001101001000001010011100110100001;
        12'd3208: TDATA = 50'b10011001011001010111101111000001010001101001011111;
        12'd3209: TDATA = 50'b10011001010111110101110111000001001111101100100011;
        12'd3210: TDATA = 50'b10011001010110010011111111000001001101101111101010;
        12'd3211: TDATA = 50'b10011001010100110010001001000001001011110010111000;
        12'd3212: TDATA = 50'b10011001010011010000011011000001001001110110001111;
        12'd3213: TDATA = 50'b10011001010001101110101111000001000111111001101101;
        12'd3214: TDATA = 50'b10011001010000001101000011000001000101111101001101;
        12'd3215: TDATA = 50'b10011001001110101011011001000001000100000000110100;
        12'd3216: TDATA = 50'b10011001001101001001110111000001000010000100100101;
        12'd3217: TDATA = 50'b10011001001011101000010111000001000000001000011100;
        12'd3218: TDATA = 50'b10011001001010000110110111000000111110001100010101;
        12'd3219: TDATA = 50'b10011001001000100101011101000000111100010000011001;
        12'd3220: TDATA = 50'b10011001000111000100000011000000111010010100011111;
        12'd3221: TDATA = 50'b10011001000101100010101011000000111000011000101011;
        12'd3222: TDATA = 50'b10011001000100000001010111000000110110011100111110;
        12'd3223: TDATA = 50'b10011001000010100000001001000000110100100001011010;
        12'd3224: TDATA = 50'b10011001000000111110111011000000110010100101111010;
        12'd3225: TDATA = 50'b10011000111111011101101011000000110000101010010111;
        12'd3226: TDATA = 50'b10011000111101111100101011000000101110101111001110;
        12'd3227: TDATA = 50'b10011000111100011011100111000000101100110100000000;
        12'd3228: TDATA = 50'b10011000111010111010100001000000101010111000110101;
        12'd3229: TDATA = 50'b10011000111001011001011111000000101000111101101111;
        12'd3230: TDATA = 50'b10011000110111111000100111000000100111000010111000;
        12'd3231: TDATA = 50'b10011000110110010111110001000000100101001000000110;
        12'd3232: TDATA = 50'b10011000110100110110110111000000100011001101010100;
        12'd3233: TDATA = 50'b10011000110011010110000101000000100001010010101011;
        12'd3234: TDATA = 50'b10011000110001110101010101000000011111011000001001;
        12'd3235: TDATA = 50'b10011000110000010100100111000000011101011101101100;
        12'd3236: TDATA = 50'b10011000101110110011111011000000011011100011010011;
        12'd3237: TDATA = 50'b10011000101101010011010011000000011001101001000011;
        12'd3238: TDATA = 50'b10011000101011110010101101000000010111101110110101;
        12'd3239: TDATA = 50'b10011000101010010010001011000000010101110100110010;
        12'd3240: TDATA = 50'b10011000101000110001110001000000010011111010111001;
        12'd3241: TDATA = 50'b10011000100111010001001111000000010010000000111010;
        12'd3242: TDATA = 50'b10011000100101110000110101000000010000000111000110;
        12'd3243: TDATA = 50'b10011000100100010000011111000000001110001101011011;
        12'd3244: TDATA = 50'b10011000100010110000001011000000001100010011110011;
        12'd3245: TDATA = 50'b10011000100001001111111111000000001010011010011000;
        12'd3246: TDATA = 50'b10011000011111101111101101000000001000100000111001;
        12'd3247: TDATA = 50'b10011000011110001111100011000000000110100111100111;
        12'd3248: TDATA = 50'b10011000011100101111011011000000000100101110011000;
        12'd3249: TDATA = 50'b10011000011011001111010101000000000010110101001110;
        12'd3250: TDATA = 50'b10011000011001101111010001000000000000111100001011;
        12'd3251: TDATA = 50'b10011000011000001111010000111111111111000011001110;
        12'd3252: TDATA = 50'b10011000010110101111010000111111111101001010010100;
        12'd3253: TDATA = 50'b10011000010101001111010110111111111011010001100011;
        12'd3254: TDATA = 50'b10011000010011101111100000111111111001011000111001;
        12'd3255: TDATA = 50'b10011000010010001111101000111111110111100000010000;
        12'd3256: TDATA = 50'b10011000010000101111111010111111110101100111110110;
        12'd3257: TDATA = 50'b10011000001111010000010000111111110011101111100010;
        12'd3258: TDATA = 50'b10011000001101110000100010111111110001110111001100;
        12'd3259: TDATA = 50'b10011000001100010000110110111111101111111110111101;
        12'd3260: TDATA = 50'b10011000001010110001010010111111101110000110110111;
        12'd3261: TDATA = 50'b10011000001001010001101010111111101100001110110000;
        12'd3262: TDATA = 50'b10011000000111110010001110111111101010010110111010;
        12'd3263: TDATA = 50'b10011000000110010010101110111111101000011111000011;
        12'd3264: TDATA = 50'b10011000000100110011010010111111100110100111010010;
        12'd3265: TDATA = 50'b10011000000011010011111010111111100100101111100111;
        12'd3266: TDATA = 50'b10011000000001110100100100111111100010111000000011;
        12'd3267: TDATA = 50'b10011000000000010101010000111111100001000000100100;
        12'd3268: TDATA = 50'b10010111111110110110000000111111011111001001001011;
        12'd3269: TDATA = 50'b10010111111101010110110100111111011101010001111001;
        12'd3270: TDATA = 50'b10010111111011110111100110111111011011011010101001;
        12'd3271: TDATA = 50'b10010111111010011000100010111111011001100011100110;
        12'd3272: TDATA = 50'b10010111111000111001011100111111010111101100100011;
        12'd3273: TDATA = 50'b10010111110111011010011010111111010101110101101000;
        12'd3274: TDATA = 50'b10010111110101111011010110111111010011111110101101;
        12'd3275: TDATA = 50'b10010111110100011100011100111111010010000111111111;
        12'd3276: TDATA = 50'b10010111110010111101100100111111010000010001010111;
        12'd3277: TDATA = 50'b10010111110001011110101100111111001110011010110010;
        12'd3278: TDATA = 50'b10010111101111111111111010111111001100100100010110;
        12'd3279: TDATA = 50'b10010111101110100001001000111111001010101101111100;
        12'd3280: TDATA = 50'b10010111101101000010011000111111001000110111101001;
        12'd3281: TDATA = 50'b10010111101011100011110000111111000111000001100000;
        12'd3282: TDATA = 50'b10010111101010000101000000111111000101001011010001;
        12'd3283: TDATA = 50'b10010111101000100110011110111111000011010101010011;
        12'd3284: TDATA = 50'b10010111100111000111111000111111000001011111010101;
        12'd3285: TDATA = 50'b10010111100101101001011000111110111111101001011111;
        12'd3286: TDATA = 50'b10010111100100001010111010111110111101110011110000;
        12'd3287: TDATA = 50'b10010111100010101100100000111110111011111110000111;
        12'd3288: TDATA = 50'b10010111100001001110000110111110111010001000100000;
        12'd3289: TDATA = 50'b10010111011111101111110000111110111000010011000000;
        12'd3290: TDATA = 50'b10010111011110010001011100111110110110011101100101;
        12'd3291: TDATA = 50'b10010111011100110011010000111110110100101000011000;
        12'd3292: TDATA = 50'b10010111011011010101000000111110110010110011000101;
        12'd3293: TDATA = 50'b10010111011001110110110010111110110000111101111001;
        12'd3294: TDATA = 50'b10010111011000011000101010111110101111001000110110;
        12'd3295: TDATA = 50'b10010111010110111010101010111110101101010100000001;
        12'd3296: TDATA = 50'b10010111010101011100100110111110101011011111000111;
        12'd3297: TDATA = 50'b10010111010011111110100100111110101001101010010010;
        12'd3298: TDATA = 50'b10010111010010100000101010111110100111110101101011;
        12'd3299: TDATA = 50'b10010111010001000010101100111110100110000000111111;
        12'd3300: TDATA = 50'b10010111001111100100110110111110100100001100100000;
        12'd3301: TDATA = 50'b10010111001110000111000010111110100010011000001000;
        12'd3302: TDATA = 50'b10010111001100101001010010111110100000100011110101;
        12'd3303: TDATA = 50'b10010111001011001011100010111110011110101111100100;
        12'd3304: TDATA = 50'b10010111001001101101110010111110011100111011010110;
        12'd3305: TDATA = 50'b10010111001000010000001000111110011011000111010001;
        12'd3306: TDATA = 50'b10010111000110110010100010111110011001010011010011;
        12'd3307: TDATA = 50'b10010111000101010100111010111110010111011111010111;
        12'd3308: TDATA = 50'b10010111000011110111011010111110010101101011100100;
        12'd3309: TDATA = 50'b10010111000010011001111100111110010011110111110111;
        12'd3310: TDATA = 50'b10010111000000111100100000111110010010000100010000;
        12'd3311: TDATA = 50'b10010110111111011111000010111110010000010000101000;
        12'd3312: TDATA = 50'b10010110111110000001110000111110001110011101010001;
        12'd3313: TDATA = 50'b10010110111100100100011100111110001100101001111000;
        12'd3314: TDATA = 50'b10010110111011000111000110111110001010110110100010;
        12'd3315: TDATA = 50'b10010110111001101001111000111110001001000011010101;
        12'd3316: TDATA = 50'b10010110111000001100101100111110000111010000001110;
        12'd3317: TDATA = 50'b10010110110110101111100110111110000101011101010001;
        12'd3318: TDATA = 50'b10010110110101010010011010111110000011101010001110;
        12'd3319: TDATA = 50'b10010110110011110101010110111110000001110111011001;
        12'd3320: TDATA = 50'b10010110110010011000010110111110000000000100101010;
        12'd3321: TDATA = 50'b10010110110000111011010110111101111110010001111101;
        12'd3322: TDATA = 50'b10010110101111011110100000111101111100011111011101;
        12'd3323: TDATA = 50'b10010110101110000001100110111101111010101100111100;
        12'd3324: TDATA = 50'b10010110101100100100101000111101111000111010011010;
        12'd3325: TDATA = 50'b10010110101011000111111000111101110111001000001000;
        12'd3326: TDATA = 50'b10010110101001101011000110111101110101010101111000;
        12'd3327: TDATA = 50'b10010110101000001110011000111101110011100011101111;
        12'd3328: TDATA = 50'b10010110100110110001101110111101110001110001101011;
        12'd3329: TDATA = 50'b10010110100101010101000110111101101111111111101101;
        12'd3330: TDATA = 50'b10010110100011111000011110111101101110001101110010;
        12'd3331: TDATA = 50'b10010110100010011011110110111101101100011011111000;
        12'd3332: TDATA = 50'b10010110100000111111011010111101101010101010010000;
        12'd3333: TDATA = 50'b10010110011111100010111010111101101000111000100110;
        12'd3334: TDATA = 50'b10010110011110000110011110111101100111000111000010;
        12'd3335: TDATA = 50'b10010110011100101010000010111101100101010101100000;
        12'd3336: TDATA = 50'b10010110011011001101101010111101100011100100000100;
        12'd3337: TDATA = 50'b10010110011001110001010110111101100001110010110001;
        12'd3338: TDATA = 50'b10010110011000010101000110111101100000000001100100;
        12'd3339: TDATA = 50'b10010110010110111000110110111101011110010000011010;
        12'd3340: TDATA = 50'b10010110010101011100101010111101011100011111010101;
        12'd3341: TDATA = 50'b10010110010100000000100010111101011010101110011010;
        12'd3342: TDATA = 50'b10010110010010100100011100111101011000111101100001;
        12'd3343: TDATA = 50'b10010110010001001000011010111101010111001100110010;
        12'd3344: TDATA = 50'b10010110001111101100010100111101010101011011111101;
        12'd3345: TDATA = 50'b10010110001110010000011000111101010011101011011001;
        12'd3346: TDATA = 50'b10010110001100110100011010111101010001111010110100;
        12'd3347: TDATA = 50'b10010110001011011000100010111101010000001010011000;
        12'd3348: TDATA = 50'b10010110001001111100101110111101001110011010000010;
        12'd3349: TDATA = 50'b10010110001000100000111000111101001100101001101110;
        12'd3350: TDATA = 50'b10010110000111000101000100111101001010111001011100;
        12'd3351: TDATA = 50'b10010110000101101001011000111101001001001001011000;
        12'd3352: TDATA = 50'b10010110000100001101101000111101000111011001010010;
        12'd3353: TDATA = 50'b10010110000010110010000000111101000101101001010101;
        12'd3354: TDATA = 50'b10010110000001010110011010111101000011111001011110;
        12'd3355: TDATA = 50'b10010101111111111010110100111101000010001001101010;
        12'd3356: TDATA = 50'b10010101111110011111010100111101000000011001111110;
        12'd3357: TDATA = 50'b10010101111101000011110100111100111110101010010101;
        12'd3358: TDATA = 50'b10010101111011101000010100111100111100111010101110;
        12'd3359: TDATA = 50'b10010101111010001100111010111100111011001011010001;
        12'd3360: TDATA = 50'b10010101111000110001100010111100111001011011111001;
        12'd3361: TDATA = 50'b10010101110111010110001110111100110111101100100111;
        12'd3362: TDATA = 50'b10010101110101111011000000111100110101111101011110;
        12'd3363: TDATA = 50'b10010101110100011111101010111100110100001110001101;
        12'd3364: TDATA = 50'b10010101110011000100100010111100110010011111010000;
        12'd3365: TDATA = 50'b10010101110001101001010100111100110000110000001110;
        12'd3366: TDATA = 50'b10010101110000001110001110111100101111000001011000;
        12'd3367: TDATA = 50'b10010101101110110011000110111100101101010010100010;
        12'd3368: TDATA = 50'b10010101101101011000001000111100101011100011111000;
        12'd3369: TDATA = 50'b10010101101011111101000110111100101001110101001101;
        12'd3370: TDATA = 50'b10010101101010100010000110111100101000000110100111;
        12'd3371: TDATA = 50'b10010101101001000111001110111100100110011000001011;
        12'd3372: TDATA = 50'b10010101100111101100011000111100100100101001110101;
        12'd3373: TDATA = 50'b10010101100110010001100010111100100010111011100001;
        12'd3374: TDATA = 50'b10010101100100110110101100111100100001001101001111;
        12'd3375: TDATA = 50'b10010101100011011011111100111100011111011111000110;
        12'd3376: TDATA = 50'b10010101100010000001001110111100011101110001000011;
        12'd3377: TDATA = 50'b10010101100000100110100010111100011100000011000010;
        12'd3378: TDATA = 50'b10010101011111001011111010111100011010010101001010;
        12'd3379: TDATA = 50'b10010101011101110001010100111100011000100111010101;
        12'd3380: TDATA = 50'b10010101011100010110110000111100010110111001100101;
        12'd3381: TDATA = 50'b10010101011010111100001110111100010101001011111011;
        12'd3382: TDATA = 50'b10010101011001100001110100111100010011011110011010;
        12'd3383: TDATA = 50'b10010101011000000111010110111100010001110000111000;
        12'd3384: TDATA = 50'b10010101010110101100111010111100010000000011011011;
        12'd3385: TDATA = 50'b10010101010101010010100110111100001110010110001000;
        12'd3386: TDATA = 50'b10010101010011111000010000111100001100101000110111;
        12'd3387: TDATA = 50'b10010101010010011101111110111100001010111011101011;
        12'd3388: TDATA = 50'b10010101010001000011110000111100001001001110100110;
        12'd3389: TDATA = 50'b10010101001111101001100100111100000111100001100101;
        12'd3390: TDATA = 50'b10010101001110001111011010111100000101110100101011;
        12'd3391: TDATA = 50'b10010101001100110101010010111100000100000111110011;
        12'd3392: TDATA = 50'b10010101001011011011001100111100000010011011000000;
        12'd3393: TDATA = 50'b10010101001010000001001100111100000000101110010110;
        12'd3394: TDATA = 50'b10010101001000100111001100111011111111000001101111;
        12'd3395: TDATA = 50'b10010101000111001101001100111011111101010101001010;
        12'd3396: TDATA = 50'b10010101000101110011010010111011111011101000101110;
        12'd3397: TDATA = 50'b10010101000100011001011110111011111001111100011011;
        12'd3398: TDATA = 50'b10010101000010111111100000111011111000001111111111;
        12'd3399: TDATA = 50'b10010101000001100101110010111011110110100011111000;
        12'd3400: TDATA = 50'b10010101000000001100000010111011110100110111101111;
        12'd3401: TDATA = 50'b10010100111110110010010000111011110011001011101000;
        12'd3402: TDATA = 50'b10010100111101011000100110111011110001011111101010;
        12'd3403: TDATA = 50'b10010100111011111110111110111011101111110011110010;
        12'd3404: TDATA = 50'b10010100111010100101010110111011101110000111111100;
        12'd3405: TDATA = 50'b10010100111001001011110100111011101100011100001111;
        12'd3406: TDATA = 50'b10010100110111110010010010111011101010110000100100;
        12'd3407: TDATA = 50'b10010100110110011000110110111011101001000101000011;
        12'd3408: TDATA = 50'b10010100110100111111011010111011100111011001100011;
        12'd3409: TDATA = 50'b10010100110011100110000000111011100101101110001001;
        12'd3410: TDATA = 50'b10010100110010001100101000111011100100000010110001;
        12'd3411: TDATA = 50'b10010100110000110011010010111011100010010111011111;
        12'd3412: TDATA = 50'b10010100101111011001111110111011100000101100010010;
        12'd3413: TDATA = 50'b10010100101110000000101110111011011111000001001011;
        12'd3414: TDATA = 50'b10010100101100100111011110111011011101010110000110;
        12'd3415: TDATA = 50'b10010100101011001110011000111011011011101011001110;
        12'd3416: TDATA = 50'b10010100101001110101010000111011011010000000011000;
        12'd3417: TDATA = 50'b10010100101000011100001010111011011000010101100011;
        12'd3418: TDATA = 50'b10010100100111000011001000111011010110101010111000;
        12'd3419: TDATA = 50'b10010100100101101010001000111011010101000000001111;
        12'd3420: TDATA = 50'b10010100100100010001000100111011010011010101100101;
        12'd3421: TDATA = 50'b10010100100010111000001100111011010001101011001010;
        12'd3422: TDATA = 50'b10010100100001011111010000111011010000000000101110;
        12'd3423: TDATA = 50'b10010100100000000110011000111011001110010110011000;
        12'd3424: TDATA = 50'b10010100011110101101100110111011001100101100001011;
        12'd3425: TDATA = 50'b10010100011101010100111000111011001011000010000011;
        12'd3426: TDATA = 50'b10010100011011111100000110111011001001010111111010;
        12'd3427: TDATA = 50'b10010100011010100011011010111011000111101101111010;
        12'd3428: TDATA = 50'b10010100011001001010101110111011000110000011111100;
        12'd3429: TDATA = 50'b10010100010111110010001000111011000100011010000111;
        12'd3430: TDATA = 50'b10010100010110011001100010111011000010110000010100;
        12'd3431: TDATA = 50'b10010100010101000001000010111011000001000110101010;
        12'd3432: TDATA = 50'b10010100010011101000011110111010111111011100111111;
        12'd3433: TDATA = 50'b10010100010010010000000010111010111101110011011101;
        12'd3434: TDATA = 50'b10010100010000110111101000111010111100001010000000;
        12'd3435: TDATA = 50'b10010100001111011111001110111010111010100000100101;
        12'd3436: TDATA = 50'b10010100001110000110110100111010111000110111001100;
        12'd3437: TDATA = 50'b10010100001100101110100000111010110111001101111101;
        12'd3438: TDATA = 50'b10010100001011010110001110111010110101100100110010;
        12'd3439: TDATA = 50'b10010100001001111110000000111010110011111011101110;
        12'd3440: TDATA = 50'b10010100001000100101110110111010110010010010101111;
        12'd3441: TDATA = 50'b10010100000111001101101010111010110000101001110010;
        12'd3442: TDATA = 50'b10010100000101110101100110111010101111000000111110;
        12'd3443: TDATA = 50'b10010100000100011101011110111010101101011000001000;
        12'd3444: TDATA = 50'b10010100000011000101011000111010101011101111011000;
        12'd3445: TDATA = 50'b10010100000001101101010110111010101010000110101101;
        12'd3446: TDATA = 50'b10010100000000010101011110111010101000011110001111;
        12'd3447: TDATA = 50'b10010011111110111101011110111010100110110101101100;
        12'd3448: TDATA = 50'b10010011111101100101100110111010100101001101010010;
        12'd3449: TDATA = 50'b10010011111100001101110010111010100011100101000001;
        12'd3450: TDATA = 50'b10010011111010110101111010111010100001111100101010;
        12'd3451: TDATA = 50'b10010011111001011110001010111010100000010100100001;
        12'd3452: TDATA = 50'b10010011111000000110011010111010011110101100011001;
        12'd3453: TDATA = 50'b10010011110110101110110000111010011101000100011010;
        12'd3454: TDATA = 50'b10010011110101010111000110111010011011011100011110;
        12'd3455: TDATA = 50'b10010011110011111111011100111010011001110100100011;
        12'd3456: TDATA = 50'b10010011110010100111111000111010011000001100110001;
        12'd3457: TDATA = 50'b10010011110001010000010100111010010110100101000001;
        12'd3458: TDATA = 50'b10010011101111111000110010111010010100111101010111;
        12'd3459: TDATA = 50'b10010011101110100001011000111010010011010101110101;
        12'd3460: TDATA = 50'b10010011101101001001111010111010010001101110010010;
        12'd3461: TDATA = 50'b10010011101011110010011110111010010000000110110101;
        12'd3462: TDATA = 50'b10010011101010011011000110111010001110011111011101;
        12'd3463: TDATA = 50'b10010011101001000011110010111010001100111000001010;
        12'd3464: TDATA = 50'b10010011100111101100100010111010001011010001000001;
        12'd3465: TDATA = 50'b10010011100110010101010000111010001001101001110101;
        12'd3466: TDATA = 50'b10010011100100111110000010111010001000000010110000;
        12'd3467: TDATA = 50'b10010011100011100110111000111010000110011011110011;
        12'd3468: TDATA = 50'b10010011100010001111110010111010000100110100111011;
        12'd3469: TDATA = 50'b10010011100000111000101010111010000011001110000010;
        12'd3470: TDATA = 50'b10010011011111100001100110111010000001100111010010;
        12'd3471: TDATA = 50'b10010011011110001010100110111010000000000000101000;
        12'd3472: TDATA = 50'b10010011011100110011100110111001111110011001111111;
        12'd3473: TDATA = 50'b10010011011011011100110000111001111100110011100011;
        12'd3474: TDATA = 50'b10010011011010000101110010111001111011001101000010;
        12'd3475: TDATA = 50'b10010011011000101110111000111001111001100110100110;
        12'd3476: TDATA = 50'b10010011010111011000001000111001111000000000010110;
        12'd3477: TDATA = 50'b10010011010110000001010000111001110110011010000001;
        12'd3478: TDATA = 50'b10010011010100101010100010111001110100110011111001;
        12'd3479: TDATA = 50'b10010011010011010011111000111001110011001101110110;
        12'd3480: TDATA = 50'b10010011010001111101001010111001110001100111110010;
        12'd3481: TDATA = 50'b10010011010000100110100010111001110000000001110111;
        12'd3482: TDATA = 50'b10010011001111001111111010111001101110011011111101;
        12'd3483: TDATA = 50'b10010011001101111001010010111001101100110110000101;
        12'd3484: TDATA = 50'b10010011001100100010110010111001101011010000011010;
        12'd3485: TDATA = 50'b10010011001011001100010000111001101001101010101101;
        12'd3486: TDATA = 50'b10010011001001110101110010111001101000000101000101;
        12'd3487: TDATA = 50'b10010011001000011111011000111001100110011111100111;
        12'd3488: TDATA = 50'b10010011000111001001000000111001100100111010001010;
        12'd3489: TDATA = 50'b10010011000101110010101010111001100011010100110011;
        12'd3490: TDATA = 50'b10010011000100011100010110111001100001101111100001;
        12'd3491: TDATA = 50'b10010011000011000110000100111001100000001010010001;
        12'd3492: TDATA = 50'b10010011000001101111110100111001011110100101000110;
        12'd3493: TDATA = 50'b10010011000000011001100110111001011101000000000000;
        12'd3494: TDATA = 50'b10010010111111000011100000111001011011011011000100;
        12'd3495: TDATA = 50'b10010010111101101101011000111001011001110110001001;
        12'd3496: TDATA = 50'b10010010111100010111010010111001011000010001010000;
        12'd3497: TDATA = 50'b10010010111011000001010000111001010110101100100000;
        12'd3498: TDATA = 50'b10010010111001101011010000111001010101000111110010;
        12'd3499: TDATA = 50'b10010010111000010101001100111001010011100011000011;
        12'd3500: TDATA = 50'b10010010110110111111010100111001010001111110100011;
        12'd3501: TDATA = 50'b10010010110101101001011000111001010000011010000001;
        12'd3502: TDATA = 50'b10010010110100010011100000111001001110110101100101;
        12'd3503: TDATA = 50'b10010010110010111101101100111001001101010001001110;
        12'd3504: TDATA = 50'b10010010110001100111111010111001001011101100111100;
        12'd3505: TDATA = 50'b10010010110000010010001010111001001010001000110000;
        12'd3506: TDATA = 50'b10010010101110111100011100111001001000100100100110;
        12'd3507: TDATA = 50'b10010010101101100110110010111001000111000000100100;
        12'd3508: TDATA = 50'b10010010101100010001000110111001000101011100100001;
        12'd3509: TDATA = 50'b10010010101010111011011110111001000011111000100011;
        12'd3510: TDATA = 50'b10010010101001100101111110111001000010010100110010;
        12'd3511: TDATA = 50'b10010010101000010000011000111001000000110000111011;
        12'd3512: TDATA = 50'b10010010100110111010111000111000111111001101001101;
        12'd3513: TDATA = 50'b10010010100101100101011110111000111101101001101000;
        12'd3514: TDATA = 50'b10010010100100010000000000111000111100000110000001;
        12'd3515: TDATA = 50'b10010010100010111010100110111000111010100010100000;
        12'd3516: TDATA = 50'b10010010100001100101010000111000111000111111000011;
        12'd3517: TDATA = 50'b10010010100000001111111100111000110111011011101101;
        12'd3518: TDATA = 50'b10010010011110111010101000111000110101111000011000;
        12'd3519: TDATA = 50'b10010010011101100101011010111000110100010101001011;
        12'd3520: TDATA = 50'b10010010011100010000001100111000110010110010000001;
        12'd3521: TDATA = 50'b10010010011010111011000000111000110001001110111100;
        12'd3522: TDATA = 50'b10010010011001100101111000111000101111101011111100;
        12'd3523: TDATA = 50'b10010010011000010000110000111000101110001000111110;
        12'd3524: TDATA = 50'b10010010010110111011101110111000101100100110001000;
        12'd3525: TDATA = 50'b10010010010101100110110000111000101011000011011000;
        12'd3526: TDATA = 50'b10010010010100010001101110111000101001100000100111;
        12'd3527: TDATA = 50'b10010010010010111100101110111000100111111101111010;
        12'd3528: TDATA = 50'b10010010010001100111110110111000100110011011010110;
        12'd3529: TDATA = 50'b10010010010000010011000000111000100100111000111000;
        12'd3530: TDATA = 50'b10010010001110111110000110111000100011010110011000;
        12'd3531: TDATA = 50'b10010010001101101001010100111000100001110100000000;
        12'd3532: TDATA = 50'b10010010001100010100100000111000100000010001101011;
        12'd3533: TDATA = 50'b10010010001010111111110000111000011110101111011010;
        12'd3534: TDATA = 50'b10010010001001101011000110111000011101001101010011;
        12'd3535: TDATA = 50'b10010010001000010110011010111000011011101011001010;
        12'd3536: TDATA = 50'b10010010000111000001110010111000011010001001001001;
        12'd3537: TDATA = 50'b10010010000101101101001100111000011000100111001010;
        12'd3538: TDATA = 50'b10010010000100011000101000111000010111000101010001;
        12'd3539: TDATA = 50'b10010010000011000100000110111000010101100011011100;
        12'd3540: TDATA = 50'b10010010000001101111101100111000010100000001110001;
        12'd3541: TDATA = 50'b10010010000000011011001010111000010010100000000000;
        12'd3542: TDATA = 50'b10010001111111000110110000111000010000111110011000;
        12'd3543: TDATA = 50'b10010001111101110010011000111000001111011100110101;
        12'd3544: TDATA = 50'b10010001111100011110000010111000001101111011010111;
        12'd3545: TDATA = 50'b10010001111011001001110000111000001100011001111111;
        12'd3546: TDATA = 50'b10010001111001110101011100111000001010111000100101;
        12'd3547: TDATA = 50'b10010001111000100001001010111000001001010111010000;
        12'd3548: TDATA = 50'b10010001110111001101000000111000000111110110000111;
        12'd3549: TDATA = 50'b10010001110101111000110010111000000110010100111001;
        12'd3550: TDATA = 50'b10010001110100100100101100111000000100110011111000;
        12'd3551: TDATA = 50'b10010001110011010000101000111000000011010010111011;
        12'd3552: TDATA = 50'b10010001110001111100100110111000000001110010000000;
        12'd3553: TDATA = 50'b10010001110000101000100010111000000000010001000111;
        12'd3554: TDATA = 50'b10010001101111010100100110110111111110110000010111;
        12'd3555: TDATA = 50'b10010001101110000000100110110111111101001111100101;
        12'd3556: TDATA = 50'b10010001101100101100101000110111111011101110111000;
        12'd3557: TDATA = 50'b10010001101011011000111000110111111010001110011010;
        12'd3558: TDATA = 50'b10010001101010000100111110110111111000101101110100;
        12'd3559: TDATA = 50'b10010001101000110001001010110111110111001101010111;
        12'd3560: TDATA = 50'b10010001100111011101011000110111110101101100111111;
        12'd3561: TDATA = 50'b10010001100110001001101000110111110100001100101000;
        12'd3562: TDATA = 50'b10010001100100110101111010110111110010101100010111;
        12'd3563: TDATA = 50'b10010001100011100010010010110111110001001100001111;
        12'd3564: TDATA = 50'b10010001100010001110101010110111101111101100001000;
        12'd3565: TDATA = 50'b10010001100000111011000010110111101110001100000011;
        12'd3566: TDATA = 50'b10010001011111100111011010110111101100101011111111;
        12'd3567: TDATA = 50'b10010001011110010011111010110111101011001100001000;
        12'd3568: TDATA = 50'b10010001011101000000011100110111101001101100010010;
        12'd3569: TDATA = 50'b10010001011011101100111010110111101000001100011011;
        12'd3570: TDATA = 50'b10010001011010011001100100110111100110101100110011;
        12'd3571: TDATA = 50'b10010001011001000110001010110111100101001101001001;
        12'd3572: TDATA = 50'b10010001010111110010110010110111100011101101100001;
        12'd3573: TDATA = 50'b10010001010110011111011100110111100010001101111110;
        12'd3574: TDATA = 50'b10010001010101001100001100110111100000101110100100;
        12'd3575: TDATA = 50'b10010001010011111000111100110111011111001111001100;
        12'd3576: TDATA = 50'b10010001010010100101101100110111011101101111110101;
        12'd3577: TDATA = 50'b10010001010001010010011110110111011100010000100011;
        12'd3578: TDATA = 50'b10010001001111111111011010110111011010110001011110;
        12'd3579: TDATA = 50'b10010001001110101100010100110111011001010010010110;
        12'd3580: TDATA = 50'b10010001001101011001001010110111010111110011001101;
        12'd3581: TDATA = 50'b10010001001100000110001100110111010110010100010100;
        12'd3582: TDATA = 50'b10010001001010110011001010110111010100110101011000;
        12'd3583: TDATA = 50'b10010001001001100000010000110111010011010110100101;
        12'd3584: TDATA = 50'b10010001001000001101001110110111010001110111101101;
        12'd3585: TDATA = 50'b10010001000110111010010110110111010000011001000001;
        12'd3586: TDATA = 50'b10010001000101100111011110110111001110111010010111;
        12'd3587: TDATA = 50'b10010001000100010100110000110111001101011011111001;
        12'd3588: TDATA = 50'b10010001000011000001111000110111001011111101010010;
        12'd3589: TDATA = 50'b10010001000001101111000110110111001010011110110011;
        12'd3590: TDATA = 50'b10010001000000011100011010110111001001000000011101;
        12'd3591: TDATA = 50'b10010000111111001001101110110111000111100010001001;
        12'd3592: TDATA = 50'b10010000111101110111000010110111000110000011110111;
        12'd3593: TDATA = 50'b10010000111100100100011000110111000100100101101001;
        12'd3594: TDATA = 50'b10010000111011010001110110110111000011000111100100;
        12'd3595: TDATA = 50'b10010000111001111111010000110111000001101001011110;
        12'd3596: TDATA = 50'b10010000111000101100110000110111000000001011100000;
        12'd3597: TDATA = 50'b10010000110111011010010000110110111110101101100011;
        12'd3598: TDATA = 50'b10010000110110000111110010110110111101001111101100;
        12'd3599: TDATA = 50'b10010000110100110101011000110110111011110001111001;
        12'd3600: TDATA = 50'b10010000110011100010111110110110111010010100001001;
        12'd3601: TDATA = 50'b10010000110010010000101000110110111000110110011101;
        12'd3602: TDATA = 50'b10010000110000111110010100110110110111011000110111;
        12'd3603: TDATA = 50'b10010000101111101100000000110110110101111011010010;
        12'd3604: TDATA = 50'b10010000101110011001110010110110110100011101110101;
        12'd3605: TDATA = 50'b10010000101101000111100100110110110011000000011011;
        12'd3606: TDATA = 50'b10010000101011110101011000110110110001100011000101;
        12'd3607: TDATA = 50'b10010000101010100011010000110110110000000101110101;
        12'd3608: TDATA = 50'b10010000101001010001001000110110101110101000100110;
        12'd3609: TDATA = 50'b10010000100111111111000100110110101101001011011100;
        12'd3610: TDATA = 50'b10010000100110101100111110110110101011101110010100;
        12'd3611: TDATA = 50'b10010000100101011011000010110110101010010001010111;
        12'd3612: TDATA = 50'b10010000100100001001000000110110101000110100010110;
        12'd3613: TDATA = 50'b10010000100010110111001000110110100111010111100000;
        12'd3614: TDATA = 50'b10010000100001100101001100110110100101111010101001;
        12'd3615: TDATA = 50'b10010000100000010011010110110110100100011101111010;
        12'd3616: TDATA = 50'b10010000011111000001100010110110100011000001010000;
        12'd3617: TDATA = 50'b10010000011101101111101010110110100001100100100001;
        12'd3618: TDATA = 50'b10010000011100011101111010110110100000000111111110;
        12'd3619: TDATA = 50'b10010000011011001100001010110110011110101011011100;
        12'd3620: TDATA = 50'b10010000011001111010100000110110011101001111000011;
        12'd3621: TDATA = 50'b10010000011000101000110110110110011011110010101011;
        12'd3622: TDATA = 50'b10010000010111010111001000110110011010010110010010;
        12'd3623: TDATA = 50'b10010000010110000101101000110110011000111010001000;
        12'd3624: TDATA = 50'b10010000010100110100000000110110010111011101111001;
        12'd3625: TDATA = 50'b10010000010011100010100000110110010110000001110010;
        12'd3626: TDATA = 50'b10010000010010010000111100110110010100100101101001;
        12'd3627: TDATA = 50'b10010000010000111111100100110110010011001001110000;
        12'd3628: TDATA = 50'b10010000001111101110000110110110010001101101110001;
        12'd3629: TDATA = 50'b10010000001110011100101010110110010000010001111000;
        12'd3630: TDATA = 50'b10010000001101001011010010110110001110110110000011;
        12'd3631: TDATA = 50'b10010000001011111010000000110110001101011010010111;
        12'd3632: TDATA = 50'b10010000001010101000101100110110001011111110101001;
        12'd3633: TDATA = 50'b10010000001001010111011010110110001010100011000000;
        12'd3634: TDATA = 50'b10010000001000000110001110110110001001000111011111;
        12'd3635: TDATA = 50'b10010000000110110100111110110110000111101011111101;
        12'd3636: TDATA = 50'b10010000000101100011111000110110000110010000100110;
        12'd3637: TDATA = 50'b10010000000100010010101010110110000100110101000111;
        12'd3638: TDATA = 50'b10010000000011000001100110110110000011011001110111;
        12'd3639: TDATA = 50'b10010000000001110000100100110110000001111110101001;
        12'd3640: TDATA = 50'b10010000000000011111100000110110000000100011011100;
        12'd3641: TDATA = 50'b10001111111111001110100000110101111111001000010100;
        12'd3642: TDATA = 50'b10001111111101111101100100110101111101101101010001;
        12'd3643: TDATA = 50'b10001111111100101100100110110101111100010010010000;
        12'd3644: TDATA = 50'b10001111111011011011110000110101111010110111010111;
        12'd3645: TDATA = 50'b10001111111010001010111000110101111001011100100000;
        12'd3646: TDATA = 50'b10001111111000111010001000110101111000000001110001;
        12'd3647: TDATA = 50'b10001111110111101001010000110101110110100110111101;
        12'd3648: TDATA = 50'b10001111110110011000100000110101110101001100010001;
        12'd3649: TDATA = 50'b10001111110101000111101110110101110011110001100111;
        12'd3650: TDATA = 50'b10001111110011110111000000110101110010010111000010;
        12'd3651: TDATA = 50'b10001111110010100110011000110101110000111100100101;
        12'd3652: TDATA = 50'b10001111110001010101101110110101101111100010000110;
        12'd3653: TDATA = 50'b10001111110000000101001000110101101110000111110000;
        12'd3654: TDATA = 50'b10001111101110110100100110110101101100101101011110;
        12'd3655: TDATA = 50'b10001111101101100100000010110101101011010011001011;
        12'd3656: TDATA = 50'b10001111101100010011100110110101101001111001000011;
        12'd3657: TDATA = 50'b10001111101011000011000110110101101000011110111010;
        12'd3658: TDATA = 50'b10001111101001110010101010110101100111000100110110;
        12'd3659: TDATA = 50'b10001111101000100010010010110101100101101010110110;
        12'd3660: TDATA = 50'b10001111100111010001111100110101100100010000111100;
        12'd3661: TDATA = 50'b10001111100110000001100110110101100010110111000011;
        12'd3662: TDATA = 50'b10001111100100110001010000110101100001011101001011;
        12'd3663: TDATA = 50'b10001111100011100001000000110101100000000011011100;
        12'd3664: TDATA = 50'b10001111100010010000110000110101011110101001101111;
        12'd3665: TDATA = 50'b10001111100001000000100110110101011101010000001001;
        12'd3666: TDATA = 50'b10001111011111110000011000110101011011110110100010;
        12'd3667: TDATA = 50'b10001111011110100000001110110101011010011101000000;
        12'd3668: TDATA = 50'b10001111011101010000001010110101011001000011100110;
        12'd3669: TDATA = 50'b10001111011100000000000100110101010111101010001010;
        12'd3670: TDATA = 50'b10001111011010110000000010110101010110010000110111;
        12'd3671: TDATA = 50'b10001111011001011111111110110101010100110111100010;
        12'd3672: TDATA = 50'b10001111011000010000000100110101010011011110011000;
        12'd3673: TDATA = 50'b10001111010111000000001000110101010010000101010000;
        12'd3674: TDATA = 50'b10001111010101110000010000110101010000101100001101;
        12'd3675: TDATA = 50'b10001111010100100000011000110101001111010011001011;
        12'd3676: TDATA = 50'b10001111010011010000100000110101001101111010001011;
        12'd3677: TDATA = 50'b10001111010010000000101000110101001100100001001101;
        12'd3678: TDATA = 50'b10001111010000110000111010110101001011001000011010;
        12'd3679: TDATA = 50'b10001111001111100001001110110101001001101111101100;
        12'd3680: TDATA = 50'b10001111001110010001011100110101001000010110111001;
        12'd3681: TDATA = 50'b10001111001101000001110010110101000110111110010001;
        12'd3682: TDATA = 50'b10001111001011110010001010110101000101100101101011;
        12'd3683: TDATA = 50'b10001111001010100010100000110101000100001101000110;
        12'd3684: TDATA = 50'b10001111001001010010111110110101000010110100101010;
        12'd3685: TDATA = 50'b10001111001000000011011000110101000001011100001100;
        12'd3686: TDATA = 50'b10001111000110110011111000110101000000000011110110;
        12'd3687: TDATA = 50'b10001111000101100100011000110100111110101011100001;
        12'd3688: TDATA = 50'b10001111000100010100111110110100111101010011010101;
        12'd3689: TDATA = 50'b10001111000011000101100000110100111011111011000111;
        12'd3690: TDATA = 50'b10001111000001110110000110110100111010100010111110;
        12'd3691: TDATA = 50'b10001111000000100110110000110100111001001010111010;
        12'd3692: TDATA = 50'b10001110111111010111011100110100110111110010111010;
        12'd3693: TDATA = 50'b10001110111110001000001000110100110110011010111100;
        12'd3694: TDATA = 50'b10001110111100111000111010110100110101000011000111;
        12'd3695: TDATA = 50'b10001110111011101001101000110100110011101011001111;
        12'd3696: TDATA = 50'b10001110111010011010100000110100110010010011100011;
        12'd3697: TDATA = 50'b10001110111001001011010110110100110000111011110101;
        12'd3698: TDATA = 50'b10001110110111111100001110110100101111100100001100;
        12'd3699: TDATA = 50'b10001110110110101101000110110100101110001100100101;
        12'd3700: TDATA = 50'b10001110110101011110000000110100101100110101000010;
        12'd3701: TDATA = 50'b10001110110100001110111110110100101011011101100100;
        12'd3702: TDATA = 50'b10001110110011000000000000110100101010000110001011;
        12'd3703: TDATA = 50'b10001110110001110001000000110100101000101110110100;
        12'd3704: TDATA = 50'b10001110110000100010001000110100100111010111100100;
        12'd3705: TDATA = 50'b10001110101111010011001000110100100110000000010000;
        12'd3706: TDATA = 50'b10001110101110000100010010110100100100101001000111;
        12'd3707: TDATA = 50'b10001110101100110101011010110100100011010001111100;
        12'd3708: TDATA = 50'b10001110101011100110101010110100100001111010111101;
        12'd3709: TDATA = 50'b10001110101010010111110100110100100000100011111000;
        12'd3710: TDATA = 50'b10001110101001001001000110110100011111001100111111;
        12'd3711: TDATA = 50'b10001110100111111010011010110100011101110110000111;
        12'd3712: TDATA = 50'b10001110100110101011110000110100011100011111010101;
        12'd3713: TDATA = 50'b10001110100101011101000010110100011011001000100000;
        12'd3714: TDATA = 50'b10001110100100001110011100110100011001110001110100;
        12'd3715: TDATA = 50'b10001110100010111111111000110100011000011011001100;
        12'd3716: TDATA = 50'b10001110100001110001010100110100010111000100100110;
        12'd3717: TDATA = 50'b10001110100000100010110000110100010101101110000001;
        12'd3718: TDATA = 50'b10001110011111010100010010110100010100010111100101;
        12'd3719: TDATA = 50'b10001110011110000101110100110100010011000001001010;
        12'd3720: TDATA = 50'b10001110011100110111011000110100010001101010110011;
        12'd3721: TDATA = 50'b10001110011011101001000000110100010000010100100010;
        12'd3722: TDATA = 50'b10001110011010011010101000110100001110111110010010;
        12'd3723: TDATA = 50'b10001110011001001100010000110100001101101000000011;
        12'd3724: TDATA = 50'b10001110010111111101111110110100001100010001111101;
        12'd3725: TDATA = 50'b10001110010110101111101010110100001010111011110100;
        12'd3726: TDATA = 50'b10001110010101100001100000110100001001100101111011;
        12'd3727: TDATA = 50'b10001110010100010011001110110100001000001111111001;
        12'd3728: TDATA = 50'b10001110010011000101001000110100000110111010000101;
        12'd3729: TDATA = 50'b10001110010001110110111010110100000101100100001010;
        12'd3730: TDATA = 50'b10001110010000101000110100110100000100001110011001;
        12'd3731: TDATA = 50'b10001110001111011010110000110100000010111000101101;
        12'd3732: TDATA = 50'b10001110001110001100101110110100000001100011000011;
        12'd3733: TDATA = 50'b10001110001100111110101010110100000000001101011011;
        12'd3734: TDATA = 50'b10001110001011110000101010110011111110110111110111;
        12'd3735: TDATA = 50'b10001110001010100010101110110011111101100010010111;
        12'd3736: TDATA = 50'b10001110001001010100110000110011111100001100111010;
        12'd3737: TDATA = 50'b10001110001000000110110110110011111010110111100001;
        12'd3738: TDATA = 50'b10001110000110111001000000110011111001100010001100;
        12'd3739: TDATA = 50'b10001110000101101011001000110011111000001100111010;
        12'd3740: TDATA = 50'b10001110000100011101011000110011110110110111101111;
        12'd3741: TDATA = 50'b10001110000011001111100110110011110101100010100110;
        12'd3742: TDATA = 50'b10001110000010000001111000110011110100001101100001;
        12'd3743: TDATA = 50'b10001110000000110100001010110011110010111000011110;
        12'd3744: TDATA = 50'b10001101111111100110100000110011110001100011100000;
        12'd3745: TDATA = 50'b10001101111110011000111000110011110000001110100110;
        12'd3746: TDATA = 50'b10001101111101001011010000110011101110111001101110;
        12'd3747: TDATA = 50'b10001101111011111101101010110011101101100100111010;
        12'd3748: TDATA = 50'b10001101111010110000000110110011101100010000001000;
        12'd3749: TDATA = 50'b10001101111001100010100100110011101010111011011011;
        12'd3750: TDATA = 50'b10001101111000010101000010110011101001100110101111;
        12'd3751: TDATA = 50'b10001101110111000111101000110011101000010010001111;
        12'd3752: TDATA = 50'b10001101110101111010001010110011100110111101101001;
        12'd3753: TDATA = 50'b10001101110100101100110100110011100101101001001111;
        12'd3754: TDATA = 50'b10001101110011011111011010110011100100010100110010;
        12'd3755: TDATA = 50'b10001101110010010010001000110011100011000000011110;
        12'd3756: TDATA = 50'b10001101110001000100110010110011100001101100001000;
        12'd3757: TDATA = 50'b10001101101111110111011110110011100000010111110111;
        12'd3758: TDATA = 50'b10001101101110101010001110110011011111000011101010;
        12'd3759: TDATA = 50'b10001101101101011100111110110011011101101111011111;
        12'd3760: TDATA = 50'b10001101101100001111111000110011011100011011011111;
        12'd3761: TDATA = 50'b10001101101011000010101110110011011011000111011101;
        12'd3762: TDATA = 50'b10001101101001110101100100110011011001110011011101;
        12'd3763: TDATA = 50'b10001101101000101000100010110011011000011111100111;
        12'd3764: TDATA = 50'b10001101100111011011011100110011010111001011101101;
        12'd3765: TDATA = 50'b10001101100110001110011010110011010101110111111011;
        12'd3766: TDATA = 50'b10001101100101000001011010110011010100100100001010;
        12'd3767: TDATA = 50'b10001101100011110100011100110011010011010000011110;
        12'd3768: TDATA = 50'b10001101100010100111100000110011010001111100110110;
        12'd3769: TDATA = 50'b10001101100001011010101000110011010000101001010011;
        12'd3770: TDATA = 50'b10001101100000001101110000110011001111010101110010;
        12'd3771: TDATA = 50'b10001101011111000000111000110011001110000010010010;
        12'd3772: TDATA = 50'b10001101011101110100000100110011001100101110110110;
        12'd3773: TDATA = 50'b10001101011100100111011000110011001011011011100110;
        12'd3774: TDATA = 50'b10001101011011011010100110110011001010001000010001;
        12'd3775: TDATA = 50'b10001101011010001101110100110011001000110100111101;
        12'd3776: TDATA = 50'b10001101011001000001001010110011000111100001110100;
        12'd3777: TDATA = 50'b10001101010111110100011110110011000110001110101010;
        12'd3778: TDATA = 50'b10001101010110100111110110110011000100111011100100;
        12'd3779: TDATA = 50'b10001101010101011011010000110011000011101000100011;
        12'd3780: TDATA = 50'b10001101010100001110101010110011000010010101100011;
        12'd3781: TDATA = 50'b10001101010011000010001010110011000001000010101011;
        12'd3782: TDATA = 50'b10001101010001110101101010110010111111101111110101;
        12'd3783: TDATA = 50'b10001101010000101001001010110010111110011101000000;
        12'd3784: TDATA = 50'b10001101001111011100110000110010111101001010010010;
        12'd3785: TDATA = 50'b10001101001110010000010010110010111011110111100011;
        12'd3786: TDATA = 50'b10001101001101000011111000110010111010100100111001;
        12'd3787: TDATA = 50'b10001101001011110111100010110010111001010010010011;
        12'd3788: TDATA = 50'b10001101001010101011001110110010110111111111110010;
        12'd3789: TDATA = 50'b10001101001001011110111010110010110110101101010010;
        12'd3790: TDATA = 50'b10001101001000010010101000110010110101011010110111;
        12'd3791: TDATA = 50'b10001101000111000110011010110010110100001000100001;
        12'd3792: TDATA = 50'b10001101000101111010001010110010110010110110001001;
        12'd3793: TDATA = 50'b10001101000100101110000010110010110001100011111011;
        12'd3794: TDATA = 50'b10001101000011100001110110110010110000010001101100;
        12'd3795: TDATA = 50'b10001101000010010101101110110010101110111111100010;
        12'd3796: TDATA = 50'b10001101000001001001101010110010101101101101011100;
        12'd3797: TDATA = 50'b10001100111111111101101010110010101100011011011110;
        12'd3798: TDATA = 50'b10001100111110110001100110110010101011001001011011;
        12'd3799: TDATA = 50'b10001100111101100101100110110010101001110111100000;
        12'd3800: TDATA = 50'b10001100111100011001101010110010101000100101101001;
        12'd3801: TDATA = 50'b10001100111011001101101100110010100111010011110001;
        12'd3802: TDATA = 50'b10001100111010000001110010110010100110000010000000;
        12'd3803: TDATA = 50'b10001100111000110101111010110010100100110000010001;
        12'd3804: TDATA = 50'b10001100110111101010000100110010100011011110100111;
        12'd3805: TDATA = 50'b10001100110110011110001110110010100010001100111101;
        12'd3806: TDATA = 50'b10001100110101010010011110110010100000111011011100;
        12'd3807: TDATA = 50'b10001100110100000110101110110010011111101001111100;
        12'd3808: TDATA = 50'b10001100110010111010111110110010011110011000011101;
        12'd3809: TDATA = 50'b10001100110001101111010000110010011101000111000011;
        12'd3810: TDATA = 50'b10001100110000100011100110110010011011110101101110;
        12'd3811: TDATA = 50'b10001100101111011000000000110010011010100100011101;
        12'd3812: TDATA = 50'b10001100101110001100011000110010011001010011001101;
        12'd3813: TDATA = 50'b10001100101101000000110010110010011000000001111111;
        12'd3814: TDATA = 50'b10001100101011110101010000110010010110110000111001;
        12'd3815: TDATA = 50'b10001100101010101001110000110010010101011111110100;
        12'd3816: TDATA = 50'b10001100101001011110001110110010010100001110110000;
        12'd3817: TDATA = 50'b10001100101000010010110100110010010010111101110100;
        12'd3818: TDATA = 50'b10001100100111000111010110110010010001101100110111;
        12'd3819: TDATA = 50'b10001100100101111011111010110010010000011011111110;
        12'd3820: TDATA = 50'b10001100100100110000100010110010001111001011001001;
        12'd3821: TDATA = 50'b10001100100011100101010000110010001101111010011100;
        12'd3822: TDATA = 50'b10001100100010011001111100110010001100101001101110;
        12'd3823: TDATA = 50'b10001100100001001110101010110010001011011001000100;
        12'd3824: TDATA = 50'b10001100100000000011011000110010001010001000011011;
        12'd3825: TDATA = 50'b10001100011110111000001000110010001000110111110111;
        12'd3826: TDATA = 50'b10001100011101101100111010110010000111100111010100;
        12'd3827: TDATA = 50'b10001100011100100001110100110010000110010110111100;
        12'd3828: TDATA = 50'b10001100011011010110101110110010000101000110100110;
        12'd3829: TDATA = 50'b10001100011010001011100010110010000011110110001010;
        12'd3830: TDATA = 50'b10001100011001000000011110110010000010100101111010;
        12'd3831: TDATA = 50'b10001100010111110101011100110010000001010101101010;
        12'd3832: TDATA = 50'b10001100010110101010011100110010000000000101100000;
        12'd3833: TDATA = 50'b10001100010101011111011100110001111110110101010110;
        12'd3834: TDATA = 50'b10001100010100010100011110110001111101100101010001;
        12'd3835: TDATA = 50'b10001100010011001001101000110001111100010101010100;
        12'd3836: TDATA = 50'b10001100010001111110101010110001111011000101010010;
        12'd3837: TDATA = 50'b10001100010000110011110000110001111001110101010101;
        12'd3838: TDATA = 50'b10001100001111101001000000110001111000100101100010;
        12'd3839: TDATA = 50'b10001100001110011110001000110001110111010101101010;
        12'd3840: TDATA = 50'b10001100001101010011011000110001110110000101111010;
        12'd3841: TDATA = 50'b10001100001100001000100110110001110100110110001100;
        12'd3842: TDATA = 50'b10001100001010111101111000110001110011100110100010;
        12'd3843: TDATA = 50'b10001100001001110011001010110001110010010110111001;
        12'd3844: TDATA = 50'b10001100001000101000100010110001110001000111011000;
        12'd3845: TDATA = 50'b10001100000111011101111010110001101111110111111000;
        12'd3846: TDATA = 50'b10001100000110010011010010110001101110101000011001;
        12'd3847: TDATA = 50'b10001100000101001000101110110001101101011000111111;
        12'd3848: TDATA = 50'b10001100000011111110000110110001101100001001100100;
        12'd3849: TDATA = 50'b10001100000010110011101010110001101010111010010110;
        12'd3850: TDATA = 50'b10001100000001101001001010110001101001101011000110;
        12'd3851: TDATA = 50'b10001100000000011110101100110001101000011011111000;
        12'd3852: TDATA = 50'b10001011111111010100010000110001100111001100101110;
        12'd3853: TDATA = 50'b10001011111110001001110110110001100101111101101001;
        12'd3854: TDATA = 50'b10001011111100111111011110110001100100101110100101;
        12'd3855: TDATA = 50'b10001011111011110101001000110001100011011111100110;
        12'd3856: TDATA = 50'b10001011111010101010110010110001100010010000101000;
        12'd3857: TDATA = 50'b10001011111001100000011110110001100001000001101110;
        12'd3858: TDATA = 50'b10001011111000010110001110110001011111110010111001;
        12'd3859: TDATA = 50'b10001011110111001011111110110001011110100100000101;
        12'd3860: TDATA = 50'b10001011110110000001110010110001011101010101010101;
        12'd3861: TDATA = 50'b10001011110100110111101010110001011100000110101110;
        12'd3862: TDATA = 50'b10001011110011101101100000110001011010111000000100;
        12'd3863: TDATA = 50'b10001011110010100011010110110001011001101001011100;
        12'd3864: TDATA = 50'b10001011110001011001010010110001011000011010111011;
        12'd3865: TDATA = 50'b10001011110000001111001110110001010111001100011100;
        12'd3866: TDATA = 50'b10001011101111000101001110110001010101111110000001;
        12'd3867: TDATA = 50'b10001011101101111011010000110001010100101111101011;
        12'd3868: TDATA = 50'b10001011101100110001001100110001010011100001010000;
        12'd3869: TDATA = 50'b10001011101011100111010000110001010010010010111111;
        12'd3870: TDATA = 50'b10001011101010011101011000110001010001000100110011;
        12'd3871: TDATA = 50'b10001011101001010011100000110001001111110110101000;
        12'd3872: TDATA = 50'b10001011101000001001101000110001001110101000011111;
        12'd3873: TDATA = 50'b10001011100110111111110000110001001101011010010110;
        12'd3874: TDATA = 50'b10001011100101110110000010110001001100001100011001;
        12'd3875: TDATA = 50'b10001011100100101100010000110001001010111110011010;
        12'd3876: TDATA = 50'b10001011100011100010100000110001001001110000011111;
        12'd3877: TDATA = 50'b10001011100010011000110010110001001000100010100101;
        12'd3878: TDATA = 50'b10001011100001001111000110110001000111010100110000;
        12'd3879: TDATA = 50'b10001011100000000101100000110001000110000111000011;
        12'd3880: TDATA = 50'b10001011011110111011110000110001000100111001001101;
        12'd3881: TDATA = 50'b10001011011101110010001110110001000011101011100101;
        12'd3882: TDATA = 50'b10001011011100101000101000110001000010011101111011;
        12'd3883: TDATA = 50'b10001011011011011111001000110001000001010000011001;
        12'd3884: TDATA = 50'b10001011011010010101100010110001000000000010110010;
        12'd3885: TDATA = 50'b10001011011001001100001000110000111110110101011001;
        12'd3886: TDATA = 50'b10001011011000000010101000110000111101100111111011;
        12'd3887: TDATA = 50'b10001011010110111001001110110000111100011010100100;
        12'd3888: TDATA = 50'b10001011010101101111110100110000111011001101001111;
        12'd3889: TDATA = 50'b10001011010100100110011010110000111001111111111011;
        12'd3890: TDATA = 50'b10001011010011011101000110110000111000110010101110;
        12'd3891: TDATA = 50'b10001011010010010011101110110000110111100101100000;
        12'd3892: TDATA = 50'b10001011010001001010100000110000110110011000011101;
        12'd3893: TDATA = 50'b10001011010000000001001010110000110101001011010001;
        12'd3894: TDATA = 50'b10001011001110110111111100110000110011111110010000;
        12'd3895: TDATA = 50'b10001011001101101110110000110000110010110001010011;
        12'd3896: TDATA = 50'b10001011001100100101101000110000110001100100011011;
        12'd3897: TDATA = 50'b10001011001011011100011110110000110000010111100001;
        12'd3898: TDATA = 50'b10001011001010010011010110110000101111001010101011;
        12'd3899: TDATA = 50'b10001011001001001010010000110000101101111101111010;
        12'd3900: TDATA = 50'b10001011001000000001001100110000101100110001001001;
        12'd3901: TDATA = 50'b10001011000110111000000110110000101011100100011011;
        12'd3902: TDATA = 50'b10001011000101101111001010110000101010010111110111;
        12'd3903: TDATA = 50'b10001011000100100110001000110000101001001011001110;
        12'd3904: TDATA = 50'b10001011000011011101010000110000100111111110101111;
        12'd3905: TDATA = 50'b10001011000010010100010000110000100110110010001100;
        12'd3906: TDATA = 50'b10001011000001001011011010110000100101100101110011;
        12'd3907: TDATA = 50'b10001011000000000010100010110000100100011001011000;
        12'd3908: TDATA = 50'b10001010111110111001101100110000100011001101000010;
        12'd3909: TDATA = 50'b10001010111101110000110110110000100010000000101101;
        12'd3910: TDATA = 50'b10001010111100101000000110110000100000110100011111;
        12'd3911: TDATA = 50'b10001010111011011111010110110000011111101000010011;
        12'd3912: TDATA = 50'b10001010111010010110100110110000011110011100001000;
        12'd3913: TDATA = 50'b10001010111001001101111000110000011101010000000010;
        12'd3914: TDATA = 50'b10001010111000000101001110110000011100000011111111;
        12'd3915: TDATA = 50'b10001010110110111100101000110000011010111000000001;
        12'd3916: TDATA = 50'b10001010110101110011111110110000011001101100000010;
        12'd3917: TDATA = 50'b10001010110100101011010110110000011000100000000110;
        12'd3918: TDATA = 50'b10001010110011100010110010110000010111010100001111;
        12'd3919: TDATA = 50'b10001010110010011010010010110000010110001000011101;
        12'd3920: TDATA = 50'b10001010110001010001110100110000010100111100101111;
        12'd3921: TDATA = 50'b10001010110000001001010010110000010011110000111110;
        12'd3922: TDATA = 50'b10001010101111000000111000110000010010100101010110;
        12'd3923: TDATA = 50'b10001010101101111000011010110000010001011001101011;
        12'd3924: TDATA = 50'b10001010101100110000000010110000010000001110001000;
        12'd3925: TDATA = 50'b10001010101011100111101010110000001111000010100110;
        12'd3926: TDATA = 50'b10001010101010011111011000110000001101110111001100;
        12'd3927: TDATA = 50'b10001010101001010111000010110000001100101011110000;
        12'd3928: TDATA = 50'b10001010101000001110110000110000001011100000011000;
        12'd3929: TDATA = 50'b10001010100111000110011110110000001010010101000001;
        12'd3930: TDATA = 50'b10001010100101111110010000110000001001001001101111;
        12'd3931: TDATA = 50'b10001010100100110110000100110000000111111110100001;
        12'd3932: TDATA = 50'b10001010100011101101111010110000000110110011011000;
        12'd3933: TDATA = 50'b10001010100010100101101110110000000101101000001100;
        12'd3934: TDATA = 50'b10001010100001011101101000110000000100011101001000;
        12'd3935: TDATA = 50'b10001010100000010101100010110000000011010010000101;
        12'd3936: TDATA = 50'b10001010011111001101100010110000000010000111001010;
        12'd3937: TDATA = 50'b10001010011110000101011010110000000000111100000111;
        12'd3938: TDATA = 50'b10001010011100111101010110101111111111110001001011;
        12'd3939: TDATA = 50'b10001010011011110101100000101111111110100110011100;
        12'd3940: TDATA = 50'b10001010011010101101100000101111111101011011100110;
        12'd3941: TDATA = 50'b10001010011001100101100110101111111100010000110111;
        12'd3942: TDATA = 50'b10001010011000011101101000101111111011000110000110;
        12'd3943: TDATA = 50'b10001010010111010101111000101111111001111011100011;
        12'd3944: TDATA = 50'b10001010010110001101111110101111111000110000110111;
        12'd3945: TDATA = 50'b10001010010101000110001010101111110111100110010011;
        12'd3946: TDATA = 50'b10001010010011111110010110101111110110011011110001;
        12'd3947: TDATA = 50'b10001010010010110110101000101111110101010001010101;
        12'd3948: TDATA = 50'b10001010010001101110110110101111110100000110111000;
        12'd3949: TDATA = 50'b10001010010000100111001000101111110010111100011111;
        12'd3950: TDATA = 50'b10001010001111011111011110101111110001110010001011;
        12'd3951: TDATA = 50'b10001010001110010111110110101111110000100111111011;
        12'd3952: TDATA = 50'b10001010001101010000001110101111101111011101101100;
        12'd3953: TDATA = 50'b10001010001100001000100110101111101110010011011110;
        12'd3954: TDATA = 50'b10001010001011000000111110101111101101001001010001;
        12'd3955: TDATA = 50'b10001010001001111001011110101111101011111111001111;
        12'd3956: TDATA = 50'b10001010001000110001111010101111101010110101001000;
        12'd3957: TDATA = 50'b10001010000111101010011110101111101001101011001011;
        12'd3958: TDATA = 50'b10001010000110100011000010101111101000100001010000;
        12'd3959: TDATA = 50'b10001010000101011011100110101111100111010111010110;
        12'd3960: TDATA = 50'b10001010000100010100001010101111100110001101011101;
        12'd3961: TDATA = 50'b10001010000011001100110000101111100101000011101000;
        12'd3962: TDATA = 50'b10001010000010000101011010101111100011111001111000;
        12'd3963: TDATA = 50'b10001010000000111110000010101111100010110000000101;
        12'd3964: TDATA = 50'b10001001111111110110101110101111100001100110011010;
        12'd3965: TDATA = 50'b10001001111110101111011110101111100000011100110100;
        12'd3966: TDATA = 50'b10001001111101101000001110101111011111010011001110;
        12'd3967: TDATA = 50'b10001001111100100000111110101111011110001001101010;
        12'd3968: TDATA = 50'b10001001111011011001111000101111011101000000010000;
        12'd3969: TDATA = 50'b10001001111010010010101110101111011011110110110100;
        12'd3970: TDATA = 50'b10001001111001001011100100101111011010101101011010;
        12'd3971: TDATA = 50'b10001001111000000100011010101111011001100100000000;
        12'd3972: TDATA = 50'b10001001110110111101011000101111011000011010110010;
        12'd3973: TDATA = 50'b10001001110101110110010010101111010111010001011110;
        12'd3974: TDATA = 50'b10001001110100101111010000101111010110001000010001;
        12'd3975: TDATA = 50'b10001001110011101000010010101111010100111111001001;
        12'd3976: TDATA = 50'b10001001110010100001001110101111010011110101111100;
        12'd3977: TDATA = 50'b10001001110001011010010100101111010010101100111001;
        12'd3978: TDATA = 50'b10001001110000010011011000101111010001100011110111;
        12'd3979: TDATA = 50'b10001001101111001100100000101111010000011010111010;
        12'd3980: TDATA = 50'b10001001101110000101101000101111001111010001111110;
        12'd3981: TDATA = 50'b10001001101100111110110000101111001110001001000011;
        12'd3982: TDATA = 50'b10001001101011110111111100101111001101000000001100;
        12'd3983: TDATA = 50'b10001001101010110001010000101111001011110111011111;
        12'd3984: TDATA = 50'b10001001101001101010011010101111001010101110101011;
        12'd3985: TDATA = 50'b10001001101000100011101000101111001001100101111011;
        12'd3986: TDATA = 50'b10001001100111011101000000101111001000011101010101;
        12'd3987: TDATA = 50'b10001001100110010110010000101111000111010100101010;
        12'd3988: TDATA = 50'b10001001100101001111101000101111000110001100000111;
        12'd3989: TDATA = 50'b10001001100100001000111110101111000101000011100101;
        12'd3990: TDATA = 50'b10001001100011000010010110101111000011111011000011;
        12'd3991: TDATA = 50'b10001001100001111011110010101111000010110010101010;
        12'd3992: TDATA = 50'b10001001100000110101010000101111000001101010010001;
        12'd3993: TDATA = 50'b10001001011111101110110000101111000000100001111101;
        12'd3994: TDATA = 50'b10001001011110101000010000101110111111011001101001;
        12'd3995: TDATA = 50'b10001001011101100001110000101110111110010001010111;
        12'd3996: TDATA = 50'b10001001011100011011010010101110111101001001001001;
        12'd3997: TDATA = 50'b10001001011011010100111000101110111100000001000000;
        12'd3998: TDATA = 50'b10001001011010001110011110101110111010111000110111;
        12'd3999: TDATA = 50'b10001001011001001000001000101110111001110000110011;
        12'd4000: TDATA = 50'b10001001011000000001110000101110111000101000110000;
        12'd4001: TDATA = 50'b10001001010110111011011010101110110111100000101110;
        12'd4002: TDATA = 50'b10001001010101110101001100101110110110011000110111;
        12'd4003: TDATA = 50'b10001001010100101110111000101110110101010000111010;
        12'd4004: TDATA = 50'b10001001010011101000101010101110110100001001000101;
        12'd4005: TDATA = 50'b10001001010010100010011100101110110011000001010001;
        12'd4006: TDATA = 50'b10001001010001011100010000101110110001111001100001;
        12'd4007: TDATA = 50'b10001001010000010110001000101110110000110001110101;
        12'd4008: TDATA = 50'b10001001001111010000000000101110101111101010001011;
        12'd4009: TDATA = 50'b10001001001110001001111000101110101110100010100001;
        12'd4010: TDATA = 50'b10001001001101000011110100101110101101011010111100;
        12'd4011: TDATA = 50'b10001001001011111101101110101110101100010011011000;
        12'd4012: TDATA = 50'b10001001001010110111110010101110101011001011111110;
        12'd4013: TDATA = 50'b10001001001001110001110000101110101010000100100000;
        12'd4014: TDATA = 50'b10001001001000101011101110101110101000111101000010;
        12'd4015: TDATA = 50'b10001001000111100101110110101110100111110101101111;
        12'd4016: TDATA = 50'b10001001000110011111110110101110100110101110010111;
        12'd4017: TDATA = 50'b10001001000101011010000000101110100101100111001001;
        12'd4018: TDATA = 50'b10001001000100010100001010101110100100011111111100;
        12'd4019: TDATA = 50'b10001001000011001110010010101110100011011000101101;
        12'd4020: TDATA = 50'b10001001000010001000011100101110100010010001100011;
        12'd4021: TDATA = 50'b10001001000001000010101100101110100001001010011111;
        12'd4022: TDATA = 50'b10001000111111111100111100101110100000000011011101;
        12'd4023: TDATA = 50'b10001000111110110111001100101110011110111100011100;
        12'd4024: TDATA = 50'b10001000111101110001011110101110011101110101011111;
        12'd4025: TDATA = 50'b10001000111100101011110010101110011100101110100100;
        12'd4026: TDATA = 50'b10001000111011100110001000101110011011100111101100;
        12'd4027: TDATA = 50'b10001000111010100000011110101110011010100000110110;
        12'd4028: TDATA = 50'b10001000111001011010110110101110011001011010000100;
        12'd4029: TDATA = 50'b10001000111000010101010010101110011000010011010110;
        12'd4030: TDATA = 50'b10001000110111001111101110101110010111001100101001;
        12'd4031: TDATA = 50'b10001000110110001010001110101110010110000110000000;
        12'd4032: TDATA = 50'b10001000110101000100110000101110010100111111011011;
        12'd4033: TDATA = 50'b10001000110011111111001110101110010011111000110101;
        12'd4034: TDATA = 50'b10001000110010111001110100101110010010110010010110;
        12'd4035: TDATA = 50'b10001000110001110100010110101110010001101011110100;
        12'd4036: TDATA = 50'b10001000110000101110111010101110010000100101010111;
        12'd4037: TDATA = 50'b10001000101111101001100010101110001111011110111110;
        12'd4038: TDATA = 50'b10001000101110100100010000101110001110011000101101;
        12'd4039: TDATA = 50'b10001000101101011110111000101110001101010010010110;
        12'd4040: TDATA = 50'b10001000101100011001100110101110001100001100000111;
        12'd4041: TDATA = 50'b10001000101011010100010010101110001011000101110101;
        12'd4042: TDATA = 50'b10001000101010001111001000101110001001111111110001;
        12'd4043: TDATA = 50'b10001000101001001001110110101110001000111001100101;
        12'd4044: TDATA = 50'b10001000101000000100101010101110000111110011100000;
        12'd4045: TDATA = 50'b10001000100110111111011110101110000110101101011100;
        12'd4046: TDATA = 50'b10001000100101111010011000101110000101100111100000;
        12'd4047: TDATA = 50'b10001000100100110101010000101110000100100001100001;
        12'd4048: TDATA = 50'b10001000100011110000000110101110000011011011100100;
        12'd4049: TDATA = 50'b10001000100010101011000100101110000010010101101101;
        12'd4050: TDATA = 50'b10001000100001100110000100101110000001001111111011;
        12'd4051: TDATA = 50'b10001000100000100001000000101110000000001010000111;
        12'd4052: TDATA = 50'b10001000011111011100000000101101111111000100010111;
        12'd4053: TDATA = 50'b10001000011110010111000100101101111101111110101011;
        12'd4054: TDATA = 50'b10001000011101010010000110101101111100111001000001;
        12'd4055: TDATA = 50'b10001000011100001101010000101101111011110011011101;
        12'd4056: TDATA = 50'b10001000011011001000010110101101111010101101110111;
        12'd4057: TDATA = 50'b10001000011010000011011000101101111001101000010000;
        12'd4058: TDATA = 50'b10001000011000111110101000101101111000100010110110;
        12'd4059: TDATA = 50'b10001000010111111001110000101101110111011101010111;
        12'd4060: TDATA = 50'b10001000010110110101000000101101110110010111111111;
        12'd4061: TDATA = 50'b10001000010101110000010010101101110101010010101011;
        12'd4062: TDATA = 50'b10001000010100101011100000101101110100001101010101;
        12'd4063: TDATA = 50'b10001000010011100110110010101101110011001000000011;
        12'd4064: TDATA = 50'b10001000010010100010001000101101110010000010110110;
        12'd4065: TDATA = 50'b10001000010001011101100000101101110000111101101100;
        12'd4066: TDATA = 50'b10001000010000011000110010101101101111111000011110;
        12'd4067: TDATA = 50'b10001000001111010100010000101101101110110011011100;
        12'd4068: TDATA = 50'b10001000001110001111101000101101101101101110010110;
        12'd4069: TDATA = 50'b10001000001101001011000110101101101100101001010111;
        12'd4070: TDATA = 50'b10001000001100000110100000101101101011100100010110;
        12'd4071: TDATA = 50'b10001000001011000010000010101101101010011111011100;
        12'd4072: TDATA = 50'b10001000001001111101100010101101101001011010100011;
        12'd4073: TDATA = 50'b10001000001000111001000110101101101000010101101110;
        12'd4074: TDATA = 50'b10001000000111110100101010101101100111010000111011;
        12'd4075: TDATA = 50'b10001000000110110000001110101101100110001100001000;
        12'd4076: TDATA = 50'b10001000000101101011111000101101100101000111011101;
        12'd4077: TDATA = 50'b10001000000100100111100000101101100100000010101111;
        12'd4078: TDATA = 50'b10001000000011100011001010101101100010111110000110;
        12'd4079: TDATA = 50'b10001000000010011110110110101101100001111001100001;
        12'd4080: TDATA = 50'b10001000000001011010100100101101100000110100111101;
        12'd4081: TDATA = 50'b10001000000000010110010100101101011111110000011101;
        12'd4082: TDATA = 50'b10000111111111010010000100101101011110101011111110;
        12'd4083: TDATA = 50'b10000111111110001101110110101101011101100111100011;
        12'd4084: TDATA = 50'b10000111111101001001110000101101011100100011001111;
        12'd4085: TDATA = 50'b10000111111100000101100110101101011011011110111001;
        12'd4086: TDATA = 50'b10000111111011000001011100101101011010011010100101;
        12'd4087: TDATA = 50'b10000111111001111101010010101101011001010110010001;
        12'd4088: TDATA = 50'b10000111111000111001010000101101011000010010000111;
        12'd4089: TDATA = 50'b10000111110111110101001010101101010111001101111001;
        12'd4090: TDATA = 50'b10000111110110110001001000101101010110001001110010;
        12'd4091: TDATA = 50'b10000111110101101101001010101101010101000101101110;
        12'd4092: TDATA = 50'b10000111110100101001000110101101010100000001100110;
        12'd4093: TDATA = 50'b10000111110011100101001100101101010010111101101000;
        12'd4094: TDATA = 50'b10000111110010100001010000101101010001111001101011;
        12'd4095: TDATA = 50'b10000111110001011101011000101101010000110101110010;

	endcase
    end
    endfunction

    wire [49:0] tdata;
    assign tdata = TDATA(index);

    wire [24:0] thalf_x0;
    wire [24:0] half_x03;
    assign thalf_x0 = tdata[49:25];
    assign half_x03 = tdata[24:0];

    wire [48:0] half_ax03;
    assign half_ax03 = {1'b1,mx} * half_x03;

    wire [24:0] mrb;
    assign mrb = {1'b0,half_ax03[48:25]};

    wire [24:0] mra;
    assign mra = thalf_x0 - mrb;

    wire [22:0] mr;
    assign mr = mra[22:0];

    wire [47:0] mya;
    assign mya = {1'b1,mr} * {1'b1,mx};

    wire [7:0] ey;
    wire [22:0] my;
    assign ey = (ex == 0) ? 0: (8'd63 + {1'b0,ex[7:1]} + odd_flag + (x[23:0] == {1'b0,{23{1'b1}}}));
    assign my = (mya[47:47]) ? mya[46:24]: mya[45:23];

    assign y = {1'b0,ey,my};

endmodule
